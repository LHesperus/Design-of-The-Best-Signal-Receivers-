��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G0��@h ���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�[@�qR�� ����"C��dKBE7\F���r����&$9g8�M>PFWD#�z":���ӳ��_}��0w�\��8׋�������N���?��m��+�ڔ�wV��?��N��j�~v��QU���T���딣0&_���X0���2|	p��rw@	@us�犱t��M,�ii^sZ��yq�`݊�|���"rG�
���}�\�.�DV	��dU�;�\����vg������W�aeYgA���z�Ś��
��H,7f�t�뾌��ߞ�:��L���om�Q*���T�KF���E�������p<�������,�\gE�y�7����򘅉��G����a�����(�I�?g�f��m����bi�ī*����b�N<��;���u��w)�SU��T�d�ǽ�*1�8�'�?�瑮��plJ�Й�m��8��r���t��U+�v��d���	u\��a(�m�Q� Q١Ӿ�$r�O��C��0�� �b�F���r�x!ڜg���p�+�8O �L#\6Į�E�=�&��D�[���(��h��CV�#3��?	M��y\XFs���RL�a)��N���m��~篟|�<�Pp�#R�S�y6�'
8�:r&@d�'1DK�5�#��ʐ�/�?�#}�{�
��R/�#3��j�f�ɨVu��7���	x]���~ВnK�k���p�C���|��X��0��F@�4%�
�V[���@��p��ʞC�ݢ�ep�O��"Hz��"��L�&Tj�P�6
� �AH��J���_a�M��RwM��;���`�(��h��$�~�MUs �~�q� \���T��U	�1�_u���V����*o��֢v��͒�&z��T�`�D�1�~�G(�����Pm�!=�y����h�}cg�I��O5 �Z��[H���1�<'"doB;sѱE�%2�}���3$�" ����f����m�!=�y����h�}m�#m��9�@���E�s-q��u���;��l)P�u��F"lܵ^�ZK�1Y6�k�8���҆�|n��q�ghY�_�X����J��Y���S>�m؆\�����d��.JKF�X��b��x
� �AH�O~=�̯�FZk ��U8�}�=n��vs!��~�MUs �̢���2���V��m[=��slc�/�<�M��}�������|���=�(��/A����;���m�!=�y����h�}M���_oH]���϶	����ę�u���;�'�� +��b)A�w�yJ�x;�������Np�,�n4_�����e68O�_��u��RL�a)P���6z�D�~篟|�sA�)#iZ&����8�:r&@P`��dpfVpb��#`^���w`q����u_��f0� ����-�l��c��=nB1�>�稅��m�!=�y����h�}�#�?�G7�Kq7a�Q`��̇����u���;���#x�d�f
�,�;�NO`�!%�qQ>B�~�e���rz�� )Te(�X��m�!=�y����h�}�G���Aj�}�aaï)ZE,�j�u���;�;N��;�Dnɴ7�x�r*�6��Ś�¢d���9��Q�Dd�(����6���e�V�-(�¦�����W�ү���u��w)�S��X3�����@��."=��	+;�'d$%MJ�Й�m�X�LGA��7�_���4�l��<u.�fa�Lm�>M�pʢ���dI״Ψ�w�Ua�[���,dԌJ�-Jdj�.n�
����k�8���҆�|n����:Vx�p*u��Uk�4�~���J�Й�m�T�#Ȃ׬��;�Ӏטw"iw4�q�M�4	�Y�����\�4�sƐ�hd	��Zk ��US����HU�6율��'�~�MUs ��y�Zk�Ž��=v �'	�?��["nq���z���J�鏈wƠ��ҿe���n �����SK���B c��(�U����	x]�<��O~���J�ޔ9����IOZ'����Oh56{�I"�c�q�CP�ba�(�N?0{l��wx0�<�·�
f��o V��	��y����/���RL�a)�G{�<�����G�/9@rk��O���@��<��7C��HM|C`r�3<0��:�.u��w)�S�3k:�(�-�~篟|���v���$2����E��j8�:r&@x7.ė)O:���?!Jf��`z$�X!{^d���J{")8�*I�����%̝��9=����RL�a)ѻtUWR�N	:.���n:�ƨ�Ob�N`�gը�d�7C��H.��T�c1����)zq�M�4=g���J��c�4��ic��S�O�4�B�!�6I	�Y�����\�4�sR���i1�����W)����VIW	I��?G�~�MUs +������\���T��U	�1�_u���*����	�����	����LO9� �Ŭ��2Dm�x]��.] �'9�����L.��6�H�.���2/�f��=V"N�^{")8�*I�ց��6 �����Y<�zd諒~����L.��6+Q)?^R7D�y�B.h�hC���(:�J�5`xt��R�m�!=�y����h�}�N�5�%����b�:q�7�<^}o?�M��;]A����@����P�����?��� �S��aY�@�Nq"Jc�l�!Hr�O��C��0��$�>��wަ����2�"�9����u���;�'�� +��v�ӫ�!NX�B���")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�;��i΀�cS���?@S:ӓ��|Q��&�N���.����'V��[��|D멼����@�Z����W�<����tТ���J/g���p��
���*,f$�7Q0- ��Ck�fÜ�2/���}����сsU%���n��/���Û�E�tw:g+��T��d^��_|��3g�ݜ��s8[Z�`
5��*�z�������D���J7"~����dY�y��
r�)�Y¹w����i��T!^z[��K�j��c���c�W_QL�ѬL�1m��+Y#_WӇ�s8[ZΑ� �}E+���c�W_QL#�̔"v��ƒ)?˳ea�8����]��
��rE���ƪϤ�Yk"1/Y#_Wӆ�q�©����0�w�)�-E����}����E���ƪϤ�Yk"1/Y#_Wӆ�q�©���H��JnXe�+�Uz�QLi/-�#�~09h�i�k1i�f1?�e�Bw�M�?_W�\I���A#|��[�m���w��L�����'�@���,������0�ea�8���
ae���K�������0��r2�􉢔�S����ީ���L�FZ�1ǝ?nQO��B�E����F}�=Ll�����,۽��8֩]=$���GZ>.�0������i� ���3�ҺIÙ=�HR��=��%ct�:��RE��]n��"�,�>E����\�vņ�Q�]�ޔiyV�[R�^Ƒ��!�`�(i3%Ah�%4
>��XP��Ȩ�wl��h�U����z~�B�wj$g"�,�>E����\�v�)��+�}��]�.�b�;װ?�p��U��֜��3%Ah�%4
>��XP����s� ]� �GR��shbvk~�#x��܃Ae��'n�^0o`�U+�PAs ����
D�ZLN�	��!�`�(i3�b9���P9b��8֩]=$�?�R��nv���N�� ���3�ҺIÙ=�HF���m¡h�5,Wluϛ�?ud��������\�v�T?�7G|`��XK���Π��yGb������l0��F��j �i7�sp>s���=1�;5��X)�z.�]�\�Y%T��BP��&��J��\��;�,EfVNN�0|]<w:�!�`�(i3x�]�V��;���Ӧ��Gjh�rO-�<i���A���U��!�`�(i3x�]�V��;���Ӧ��Gjh�rO-�=|-�e1|E�A�2�����x�]�V���rژY*��5|�}KL?-���o)�]rN�ǁ�f�T�J��H9��\�v�T?�7G|`�h�May\Ƒ8P��1pri��i�����8�TP�=5Y �������w�b	�Y���S@��Q�J!�`�(i3x�]�V�� �Gk	�}���f���w�D��y.�t��rcZH���N��S�I�Q%CJHn��z��r9�3`���*1�P�9�L�,d�%$!R��!�`�(i3A( ����_ֲ��mŹ�[�g�DPp�A�h��+Fen����9��#�B�sYC��\�v��_�R�G�$����{v��G�K$xE�p4rqG7��u*K6H �i7�sp>�͹ ��I�Q4p�/�;ϔW�~p�~{H��)w�<�_N&�G"�2���k4�͹ ��qC��~�;ϔW�~p�~{H��)w�<�_N&�G"f�x��rޥ�6�DXK��]c���H������i��E����F���8�TP�}{�Z
M{2jR�j���m l�o�����!�`�(i3x�]�V��w�7qyX�񙗡��\��T}u��Q��L(\Ӧ�$�̎�)NC�lԇ�-{�v�ј�"��Z鎬���������o�	�7��r�=N�By3��<�]�!����M[��Ǣ&��s���q�����5	���]���>����C��N���u��"i��?^���-��%M�rs�i��@�N3,(��&Q��3�ց���=��"X��[����fbK7͍��|��W&":�X�=)�H�7M��񇬦���
L'���Xw��+x�r�2�6�d�f�]2�y�Z鎬����(��eظ�=�tneX N�By3��<�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e�,���6+�\.�l����"B��$I��w��,c�A�L'z��0N�7;�¬pX��g��U-�e�,���6+��kv޶Glbq�Z��T�I��w��,c�A�L'�b��9X�T��&��;�¬pX��g��U-�eaԗ5��C�6�ǌ�lA�1�:�Ω�[@�qR�� �����u���k9��0�S�&�����"m�K7{�>P�2-i_���F�� �yz��$6ea�8���
ae���K������I^wm&�BN>�4�
�����Bdʨ,��偋:�Q	Q��|��Ӻ�(,��y�ӓ������ �V�ޒ֙f���_����}�\�����Ք�)�"JHn��z�c����,XL��=d��z��_#Ԡ�T��Ɓ��~�26��\�o�mW��y�ӓ��Dc4Ƥ S!f#���������l����O	%K��ͪM$յ[+8��"Ě��	s�_�5��ǈ�A0
��_�P[f���Ն gWVbT+��uL-���S8�,������9��
����	�|���/��@���#��M&s��'�PD������Y�L�FZ�1ǝ?nQO��B�f�8
��u��r��f���ՆnZ�va�?��Ԝ�G�ǈ�A0
����m���Yk���y��j��kj�����N��U���q��m"b��_��.V��(������}Dq�f�HN��R���מu���'�N�T~�m�ڨ�hծ���%>�rGO�D mWNHN��R���מu��� �H�0��
�5ߧE4��ʥ�nr]�b�N��?�{�XԲ���:'�>����߰r�n���D�߼
�d����ň�3Of'�����4�o�r�\Tȭ�3���r�<����M��_(����@҄���G��A"�U���w�c*��t+��I���XP��Ȗ�!�Rd=��¾ȼ�����Y�L�FZ�1ǝ?nQO��B�f�8
��u��r����َ�,�f�d��j�W'� h�ҩ���=�g[V��M*�/3o�U�r*A&-�Ri����l��M�r!�B/(�B���l1tSjv�!�`�(i3
ҭ�3���O���w�_f!�`�(i3��Ě�����}Dq�f��u��A�0�Ή*��a��2S����R�5ߧE4��	��x�(�6k�4d��!��Z!�;'�F&�MB˖�4,<��Ě���z&v��\�����3�}@��9�ڮWm�pi����Q$n�ti��|�@T��޹�{kb; ����ܕ����������a�"�Z�>)��]�B���[�.��|ȃ�$����T����i-}�����&;�8��������@|������]�^��� _�HN��R���ء�I����hڻ��:��L��O��݄�$��F�Ճ����\&�}u�i��|��
��(����{��ۮ�/���YЏs/�i���M4��S�$j���f����lNȲL���"��y�X�:�.�AY�@�W���� 2�AY��)��c�H(�亠-��fn�����I�#��Zb�JHn��z�c�����<�W�C%���6V���~�26��\�o�mW���'n�^0o���˟y��èV7�%M�����$j�@��+X>N�q�p�e6�_���|(�6k�4d�{j���d��,3y�@�VҒm�fF�5.]�����������0u�\k|aT��3G���(p��1Pw�������#p��H��R��Y��[�нx*�U	s����{`F�I6��M��^P�h$;���pM���ksdDH����'n�^0oq-���N>�4�
��,���Q��b�s6�d+��#	T�d����'3��	�;�j�"�[u��C@��AO}$|~�K��������� 2��L����ֱ�q������m�q�)Ў6dG��O����14�7'U�1�R�\<۳�<�G=}Id=��¾ȼ5�����}Y��	}�@�'�C%�-"�I5]l�����zQf�H����3bQ=�3�� �֤D�A��*ȑs��-�����y��j��kj�����N����"���jVѭ@;�jmT�#z&̴T	�et�f'%<7�lv���gWw��-����!�`�(i3�zk����\��;�,�Ra])n#���r������Aڬ&W�y��v���z��N���!�`�(i3�<�I��y�G��C�m�]6^�Y�ѓ,��|��H!�`�(i3)�{6�U���Ra])n#���r�����y��j��kj�����N�
\�n/S-��}Dq�f�HN��R��bP�63Z�tHN��R���O>�R�`t�td���5��Ě����E�i�m}6�E`���ʥ�nr]�b�N���pl�4ʀ���ߦ ����Rn�pPip<ɯ�nv��2������開k����6U٤!Q
���g��Vܙ��t�cُ�Ջ6�x�p�=����w`q��La��Y�E����m�s�*�MOL�ӯ.���w7G�����]\{���bq'���7ג��W!�͘�<�W�C%���6V���~�26��\�o�mW���'n�^0o<H�-��*{y���� �!�fLf��),��9��"!<���+�37y�����:���f���,�';:ZËF�3$����Vܙ��Lߝ-�Nr��VYW\-@��F~*7���&�_],)��v@˼�\�v��\aьIR=Z�˙}���.ᬵy��Nn"��%[��o@�?� Zh�R?�R��n�#ٷ�Ef��dט�w����j����r�C�M$�&d�X0�� ���3�ҺIÙ=�H��M����A�m�(����3�y�ܓr��G(h���i�K�g;�\��f9��NJ������@zLо$ԠI�*׿j�h�<�&d�X0���E����F�'n�^0o<5������U��֜��3��P=@��������$��Xo���~��1�51	�<����ry��cTx z�Jm]A�/����<.+6J!�5����`K��� �"�W�A�&hH\!�`�(i3�b9����lY1�ËF�3$����Vܙ��|�CY�oO���^��t���9j.�l>'�o��&L���W=D��'n�^0o`�U+�PA�5����`K~����G귈nIg�R���]6���b9���P9b���dט�w�����{�������}>p~z�r,J����!_�IÙ=�HB�q;�~ =����V��g��cH�wA�?��6a/�j�m��\�vňu�,�s�p�m~|��`.t��J��|�����IW�A�&hH\l0��F��j�q	k���A�P4ǲ I�g�R����z'/)�� 0�s]7�r޸��zL͊�q��o����6J��z�h��4�*ܑe�W����n�4�c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e���b P�|h{�T��`�)�	�%{�;���;�L���9�D_�3���U_�+X���=ў@'���Xw�j�7��Vx�%L��W��_�ړ8���/�C=2崝��b�7���U��+�Xa�H(�˕�%LH�N3���XP���f�Nd+l�Yҽ֗��D)�q]�i��E��T�
���A.o�G�m�?[���S��IÙ=�H��H(�T�O��{Tɀ���S�<Ԣ�E,�J�|R�ZLN�	���P4ǲ ��V �-�{q�����/��+l0��F��j#w���	(���B��j�Q��9�V�ݦ\�t!�ǿyXAm�� ��<��]��i�"�`�|��K�z��|����=%+]Bo�A;h�F��O�i���AԢ�a\蟖�S� ?�0��E|�,°������R�wX���dט�w����j����r2��������������JHn��z�>�ack���A�;�֋`N(��/��<`�.M�� ��˽��r� B^�.�ߘ�)�I0M�/�s���'n�^0oPpkiq�o�H�MPq6.��[�#m}�
�?�A$�ʁд����-VL���+�J��Y�{'%s�O��W��-@��F~*7���&�_�EOs\�̞��>�h�5,Wlr�r%)cA�z���a�R�wX��}�
�?�A$�ʁнv1a{J�-���Ƚ�0Y�{'%s�O��W��-@��F~*7���&�_�EOs\�̞��>�h�5,Wlr�r%)cA�z���a�R�wX��}�
�?� ��U�ϴ����-VL���+�J��Y�{'%s�O��W��-@��F~*7���&�_�EOs\�̞��>�h�5,Wlr�r%)cA�z���a�R�wX��}�
�?� ��U�Ͻv1a{J�-���Ƚ�0Y�{'%s�O��W��-@��F~*7���&�_�EOs\�̞��>�h�5,Wlr�r%)cA�z���a�R�wX��}�
�?� ��U�Ͻv1a{J��8�P��Άg��dT�W/S��8(�E���Kt���pm��)|#9���b!��u�ϟ��7�4�-�`~ ��#֫��/�*ܑe�W����n�4�{lGD�V�Bf�Nd+l�Yҽ֗�6��H��q���N�t�3���_���&#ݟB�E`^n�&�
_�n�@/%{�;����f�kN�ı*�7`����\Z��K��i3�|)sՀ�/V��������A@"�,�>E��k�:A�	S�r��AR1<]Q�I����踫g(�r�N�ǁ�f�TB��vC8U�@����gG���:���U?�G%ZQl蝌b�Bϱ��ᵉ3��鑘2����.0��jOT���hLP��2�q�7s�9���o��S8�/ #O�)�����}>p~z�r,�L;Л��|#9���b!��uፂ�6J�Ko��E�`JcU#֫��/�*ܑe�W����n�4�{lGD�V�Bh�5,Wlr�r%)cAh�߆��y�����DzL�ł)w���)]���&5j�d�٣��c�A�L'�R�M`Si�c�n�R�HM���#ga(􆿳�ټ*w2�56�
�CӞD�+5�4��c�%��)� BM���1�
�]�!��	Ǹ�y85��O�\�l$�L�溥����v�8:ۛ@W:���#���F]����.Zx�.����#���Ʒ��t���(�犽{Tɀ�$����nQ�rVt.�N���G��{�ݤ!�8���/�I����"�]�N��&�|���|��] 1�0µ�]�!����w�Հ�����DzL��T�B�X
��չ�Ad��d�٣��4�5_�o0b!��u�)���A7��M�����d�٣��c�A�L'�O�({���p~z�r,���^���2������}(Q6D����d�a�4$�b!��u��V����Pјq���U��@����gG������0w��z䮃��ġC���}�
�?�`)[�-hnqo)}>�	�ғ�vq���q�41&q^�`
�c��><�$2��Я�R�wX��}�
�?�`)[�-hnhG�W�ғ�vq���q�41&q^�`
�c��><�$��;mQ��8���/����,D��ǉã1Xɟw��D�A(g
�]�*��q�41&q^�`
�c��><�$2��Я�R�wX�ո@����gG�DI߃���iA'R�	�_��<��E����FZ鎬����
C��8q��f�kN�ı��U��+�Xa�H(�˕ #EO���h{q����'6���;8=�g��U-�e,%�0g�����L���N�b�'Be�)\���!�`�(i3�[�l\�`�|��K�z��@d��ץr�&U������G|M�Y�Q��*7b!��u��N�|�c�$�t�!�`�(i3���+�J��Y�{'%s�[�&B�踫g(�r�x�y�Zgl�k�������NI�:7�N�5�%]���a(􆿳���2����.)}���/�;���_!�`�(i3!�`�(i3�􇃬Tk�H@H�֦g�㎏qló��@d��ץr�&U������G|M��=����)}���/��C�x!�H�Z���,�!�`�(i3�U,�(�)8Q�y�� Y{q����'6���;8=�g��U-�e,%�0g�����L���N�b�'Be���`F��~!�`�(i37s�9���o��S8����ٺ?�n���㬺ƃ
ᾆ�x�T�\ ��i3�|)sՀ�Oi9L�:�k]m��y�1O�r^�!�`�(i3xZ��j�
�����1��;-;*�7��;mQ��8���/����,DTc�~y��i�v1a{J�O+T-rcs�"�,�>E���]�!��	Ǹ�y85��n���F�r�f�t���ӯIJ ��`y�����g�,P�n�R<���Յ!��4�c_����+#��.X���*"v%)��Qcm hP"G�wk�P#7!smWF�r�f�t���ӯIJ ��`y����@����gG�DI߃���iA'R�	��.���E����F�R<���Յ!��4�{lGD�V�BnQ�rV��q�t7i3�|)sՀ�Oi9L�:�k]m��F���d H��(әxZ��j�
�����1��;-;*�7��;mQ��8���/����,DTc�~y��i�v1a{J���ǔ���'�P$��<�7��V�����T�=�;^�6#9���k��$a(􆿳��Y��$�	b!��u��Ɔ �����O�����PX�÷�������;^�6#9����!@�+ufw5~�.�.ᬵy�����3��
3h}Nw���85Zt�����V?�ƇBHx\�'���Xw s4S�'�i��`�z������ִG�ĵ�I7��-5��6��	���`y����@����gGI��l��i�g���:�a��Y�{'%s�[�&B�踫g(�r��C�M$�#ã�fޅ������ϲ�CyW�f�tR�wX�Ղ�hF���H#
ZM��L~΄gO�3����?��ҹ���+F�+�V��+�_��<��d�٣���������ݹ�0���f�Nd+l��p��;z���>)0'6���;8=�g��U-�e���b P�։-�.l?���݇�T%{�;���;�L���9�D_�3���U_�+X���=ў@'���Xw�j�7���d�uY�ة�;mQ��8���/����,D�I���A���]�^�kvo�Apw�I�N�_V�ܔp�l
d�R�.��On: +*��YN�ǁ�f�T���j����^��E���!��=T,��1�~�� �(׸���-��i��+b!��u፞�f
t斃����u_7s�9���on�-�6��
�jW��D���M���R'),��`��wu���뿼��8��''6���;8=�g��U-�e���b P�~?�b�e�2����t$I+�V�6IWJE�r���秹�3I^�v�[�9q�Y�{'%s��.|Z�����8��''6���;8=�g��U-�e,%�0g����A�YHm��G�m����E����F�i�_:�ܷ��	N^�U{xN��i>w��˪?�-�l~�U�n��(���(w�.#�U�EOEe�1<�6�n����=��H�Gc���=B<�O}����~�k�Q�)�v���|ۈ�٥��m��_t��:ʰ���w`qԴ�~`����vQ� ��}�
�?��,��	r�:M�'$�*��BL�Jx��e�2l��4��a��se�ξ���I��RhF���k��76�C=2崝���^�9�8pQ�J��7��!�`�(i3�Q�^�y�����9�!�`�(i3!�`�(i3!�`�(i3���Z1`�N�ǁ�f�T��	��S��H(�T�O��{Tɀ���S�<Ԣ�E,�J�|R�ZLN�	���P4ǲ �p�o*G��&1����L��h���vv���"	��� 2�I�Û[����N���gx$�O�Җ*���X�w�)?����t}�ݓ�ZeUM�ٝ�z*N�I�l�u������P4ǲ �p�o*����/�Z�k�ʆ-���t�]¥S��� 2�I�Û[����N���gx$�O�Җ*]��z�o̈�^d\�f�� l�o�bw��H(�T�O��{Tɀ�$����nQ�rV",�Ű�
iEE�G�p�o*��NB�D�u�y����R�`7�K����'3pk~��r�<Uee�N�����a"��-K8��C��Jqõ�偋:�Q	Q��|��]1B�]�b�C�r�X��À��#�P7��ŧ �GR��shbvk~�#xǩ"�4s2nQ�rV",�Ű��dט�w��^���֮�v�@[�JJ1��P�M��Ln��S�WY_���P[!�`�(i3!�`�(i3!�`�(i3"�,�>E��C.W26K�~�a�o�yai�7]����'�C}���� oI��RhF��r��,����g�,P�nv�@[�JJ혮��רc_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85�9)e�AjL�E��w*�t%��zxa(􆿳��?ƾ�s��	��6��	����}M�l8�	
ږ�|����=%+]Bo�A;h�F��O�i���AԢ�a\�W__XOhGp�&���A�]I�3Ԩg��U-�e���b PbL}b����*���G��4���r�W+`�x�of'%Th�� �GR��shbvk~�#xǩ"�4s2nQ�rV�}!�@�?0����s�Y�{'%s�O��W��W���}���i�����dq�8���/����RY��Ɛ�<["��+�O�JT��8D��V�6IWJE�\��[�B�L�溥����v�8:��|`��'J�	�LÆ��E� )�&�VR5�����b�Bϱ�r��������]�Y����f�՜�T�\ ��y�.�`L�.@E~J��g��$���M�;�E,;��0����GI$��ǂcY�~�s<��MR*����%���$������ظ@	,���:�<�L�E��w*e�΢���v��J2N��c_����+#��.X���*"v%)��Qcm hƐ�<["��+�O�/�#��P�h}Nw����x�/�c�ۡ���Z� ��(HU�î�D�p�&���A�2��:�k���`�z��Y��),�B۸��L� s�j8&��f;�P�=��X��/D$�"��! Y�]�7Syv�J�Բ�������@d��שI4��欱���j���-+��B�G}ϼ 8���hy�`�w��v1a{J��ٱc����Ɛ�<["���܁�_�0�ΩyO^~��M����A�m�([}�@��L�7�b�����x�/�c�ۡ��F</h,魰d�/�p�&���A�&�ʜ��q?H^��2踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ��{�j��<�ao����O����Ft��7G��L�E��w*e�΢���v�2��:�k���`�z��Y��),�B۸��L� s�j8&��f;�P䒡�3����me":l�n Y�]�7Syv�J�Բ�������@d��שI4��欱���j���-+��B�G}ϼ 8����n�Jt�g�v1a{J�=���c�(~Ɛ�<["���܁�_�0�ΩyO^~��M����A�m�([}�@��L}�
�?�^)�G�B�+�WdM4@��͒r��ǩb�W�[r��-�W.���g/��ξ���I��RhF���k��76�I����"��)׺������Y�U���i���@)�l��0�L�E��w*e�΢���v��J2N��{lGD�V�Bf�Nd+l�Yҽ֗��i�ܰAb!��u�zk���������XIb!�`�(i3GYs��$;���$���M�;�E,jZ"]�Vp踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ�)׺������Y�U��3Y��P4���U�L�E��w*e�p�������
��M����A�m�([}�@��L}�
�?�u����p��8��V\⯜�'�,LFb�W�[r��-�W.��@��i�=�f�kN�ı*�7`����\Z��K��4����/�Ӝ�z@����U��@at3Y��P4�\�7.��v�@[�JJ혮��ר�bl�_�p�ξ���I��RhF���k��76����,D�ʥ��G�M��K��'�,LFU�î�D�p�&���A��J2N��{lGD�V�Bf�Nd+l�Yҽ֗��i�ܰAb!��u�zk�����>�P,љI� ���۫�d�٣����Qq�M��H�_�ЩI4��欱���j���-+��B�G�
�CӞD��=2���H��̣������G���]�!��[@�zZ��g�f�kN�ı*�7`����\Z��K��4����/�Ӝ�z@����U��@atA�ᴽ��d�1�~�Z鎬�������j}�c��`�z��Y��),�B۸��L� s�j8�-D���(���!G�{s��?������H�^M'���Xw�"O=��踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ��K���B�V�C��k��38�h�3&�N�qB���'���Xw�"O=��踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ��K���B�V�C��k��38�h�3&�u�p���n�]�!��[@�zZ��g�f�kN�ı*�7`����\Z��K��4����/��)}���/����ly�P�r��n�Ŀhw�)��Ov�@[�JJ혮��ר�bl�_�p�ξ���I��RhF���k��76����,D\X��!��x�D�Re��BE�tU�î�D�p�&���A��J2N��{lGD�V�Bf�Nd+l�Yҽ֗��i�ܰAb!��u�t�,�NL}�="��x8I�3L�*}F�GYs��$;��H��,���E���:��`�z��Y��),�B۸��L� s�j8��h��)ew���m���BE�t Y�]�7Syv�J�Բ������sl����?r�<Uee�N�����H�OM��`�@����gGdR��Ƈ�r��F�f�J�v���+p���X�o�!���	����}M�l8�	
ڶ�@d��שI4��欱���j���-+��B�G3�+��m\n�v�ĺ�(���!G�{��yn_Fu�Ɛ�<["���܁�_�jZ"]�Vp踫g(�r�N�ǁ�f�TpD��ZOU����q�f@&��f;�P�=��X��/�ب����b�W�[r��-�W.��@��i�=�f�kN�ı*�7`����\Z��K��4����/��.������FD>�v��Pn<����X�o�!���	����}M�l8�	
ڶ�@d��שI4��欱���j���-+��B�G}ϼ 8���hy�`�w��v1a{J���MB��)p�&���A��J2N��{lGD�V�Bf�Nd+l�Yҽ֗��i�ܰAb!��u��@��A���k]m���r��y��L�E��w*e�p�������
��M����A�m�([}�@��L�@����gGG5������{��U����d�٣��c�A�L'G~��6�7;-;*�7��;mQ��8���/����,D�;����;�;��O�"���Q]� _�rs�i��@�N3,(�;^�6#9���k��$a(􆿳���2����.�N��+�j����tL������	�Z鎬�������(����S� ?�0��E|�,°������R�wX��}�
�?����Н���A�Y��|w�j<�lb�rs�i��@�N3,(�;^�6#9���k��$a(􆿳�P<t8��3����開�E��ч¼xE���8��w���ȟ���8�M�$�愉V�Sup�xg쬉� }���n4s1��7�癆cg3bQ=�3�� �֤D�A�f�8
�������&S��e	�/a��@�f���I4��欱���j����XN(�U�]���=�w�Ηե>���Q=z����9�r�)۬
�,#�����K1P��8?W!t��_A�;�֋`N���}J�|���|���j�)6)-
�5ߧE4��?�{�XԪ��]^)��\�׎w�-��8n$DI��'����0/ܤ�(g��V���[b�I���\�v�n��l����:%��Z��4��.�w}?�(��y(���B������P�I��RhF��K�X:��3����s�c�����gv,��u(q��Ϝ��*@&&r��]������4���8���i�_(����@҄���G��b�i0[����8|o����q,� L���,�F�?��jO���a�N����+���LQ�{p�uR�R�W�u)hZae;s9=3
���k��7)#c��Y�7#�xIQK*QYc����it	�T$x�����}�	76�&�� Ӗ�tJ��K�]���!E'�"�F�+��^�6,!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3����n�I��'����0/�e��9�S���ތ�1��\�v�n��l����:%��Z����}�%��@��I����"���_�Ps޴�ik]�7A��(�n��rs�i�� ��*b�+W���F�^�Y�7#�xI��;mQ��8���/�C=2崝�Q�gL#A=�����ׄ� a
��Vx^��\�v��|z���m��P���ݪ��*h���'�a+��tI�F�;���N%�:+W�5����`K��0)]��w�b^X�P�NI����l>o��|��>�*�).zVW�ȏ�k��a�s+�ҟ�r/�^��D途�؎���ɿJ�:9�2����rR#K�pl� �PP��ƿ�c �B�dH�7DR�i�Ρ��˧T������X�p0�&�����Q�a5���nXZjwi�U���Mչ�����Y��n�Z(Ρ����u�PBxN��X*d��Uf�Y9��_QzMy㥁�hK�'�njVfV)~�`V%'�\�*�c�E#
D�@���b~��Z��=N��!�`�(i3�d�٣��c�A�L'J����l�!�+���LQ���"X��[��Q[R�7�n~�x��<�,���E�!�`�(i3�n`5�fK�\w��0]b!��u��չ���1|���Y�ǒ��Q]� _ό���.Ӹ@����gGWm?"<��_�S�
utY�{'%s��.|Z���I7��-5��6��	���`y����@����gG�[bGf�_�S�
utY�{'%s���'����C�`�/�t�KV*�3?�|��T�5�d�,WT	W $V��8���/�I����"�nx��hѧ�F��6��U,�(�)8���0y�	 ���t��h�/a�'�̗�����C�M�����T�\ ��i3�|)sՀnx��hѧ���Nz�
���U,�(�)8���0y�	 ���t��h�/a�'�̗�����C�M�����T�\ ��i3�|)sՀg�j*8a�.F��6��U,�(�)8���0y�	��sC��#���FӪ�c�g<�g��U-�e,%�0g���p+�@�����NۥUn����n{�_�\[$Q��
�̞��>�nQ�rV�}!�@�?0a(􆿳���2����.�t��������˃�Iy��Fp����f���,(���B�����(�犽{Tɀ��k�V\���"X��[��Q[R�7kѶ���� �oi���:FI�������b�Bϱ���w�K���1`��vߜ�*�l8�b(������#oM|#9���b!��u�],��%s��O©K���AԢ�a\��F�dHB�Fvͧ"�f���-A�¤�x.�Knq�z���a�R�wX��}�
�?������3�K�?\B�]q��T�ٮ|�,
���1��e0����yN��7��aq���E���ss�T�\ ��)�g.�F�_�u��Y'G-+;X����Jn,���`ό���.�}�
�?�ʬw�S��зq8�Ј'���Xw���,DH�v������g0TF�'�]�!����w�Հ㸮�U�M��	[�/��87s�9���o��S8�l7�EL��>0�1ۍ�h �=���"X��[�d�a�4$�b!��u�V@���gx2�n`5�fK�\w��0]b!��u��4�	��`��@��⋌�U2ރ�8���/�����s�c�����gv�h�ц� )�\�~xy�Bp��!�ʆ�In��tw�?�b�>޼�\�v�	�+�&I(&�L����6�{�Pe�E"���m�PU}������[��p#ِ.��҆�3�>0�1ۍ�h �=��h��a,JD�_�k�W�A�&hH\{UY�Z�[2�h �=�)�����g�P�e�97�i��'���L�溥����v�8:hJ�tV�nQ�rV� �L_K�*��M���R��ӟ-��NiघM�.�� �i�aYB��#���Fν��E���w�w:��y��j��k[:�ۤ�U2̥�0�L�p~z�r,���Y���hvl��9�h �=��l�I�SCp~z�r,o �#^{���y����b�Ա,��H(�T�O��{Tɀ�$����J�	�LÆ�c�9ʼ��$�G�nJ `G�p�P���� ����F��O�8�c{}�C���B��	��u8-�_��C`N�r7�r��#[��Y���0�ȷS�J���4�����\�v�n��l���m�-H�h�U�p�ջ�D�T�'��k$Y��C�9I��@��F��6�!�`�(i3y��Fp����f���,(���B��\���V#��p~z�r,�b��r�
R�wX��}�
�?�oj�+p�K�J�iN�S!�`�(i3�E����FAԢ�a\��F�dH��|c_�m��ġ��,�z���a�R�wX��}�
�?�Qw�$��Z��/�dW%�!+���E����FWS���
��ʅ�-`JX-�ܶ�0l�x����b�'Be��
������n`5�fK�\w��0]b!��u�v�A�
^^3�V�C��k�HvL)���	���hF�]�!����w�Հ�JX-�ܶ�0l�x����b�'Be��
�������+NonR[�q���U��@����gGP���Ʃ8/Tu�����_&����ʺ�;[��]�!��	Ǹ�y85�A�'5�i��|�����I�HM���#ga(􆿳���2����.\�#$�ÙAWfי�b��}!D̅����<!GO#зq8�Ј'���Xw�j�7��[|��;�ċ�lʥԆ�V��,ۦ�T�\ ��i3�|)sՀ�}l�����@~H��k]m��n�_��-����Q]� _�rs�i��~�g�t�qN�c�B���)%O�lg�;S"��<[$��`y����@����gGP���Ʃ8/Tu���Ŝ��%ٿ�j;�Jw�зq8�Ј'���Xw�"O=��踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ�}l�����@~H�k����`T�]b �!�`�(i37s�9���o×��̙�F�9 }�m�f�Nd+l�Yҽ֗��i�ܰAb!��u�v�A�
^^3�V�C��k�&�c���d��b�pAзq8�Ј'���Xw�"O=��踫g(�r�N�ǁ�f�TpD��ZOUZ��| �Ɛ5�e`��9����dz����NR�p�'q�-��nEg�N>Z�k���@��b�Bϱ���w�K���1`��vߜ�*�l8�b(������l__�I����J�����g���R�wX��}�
�?�u����p�����+X��FJ���--f�`���$"�,�>E���]�!����w�Հ�b02�O�0�5G,��Gc#�T�Ed!�`�(i3��Q]� _�rs�i�M�����geE�vx���ƚP�& 5f��e�T�\ ��i3�|)sՀ�)׺����\� C&����q��Z���2%�ɛ'�F7�Gh`��@�����0y�	�l�f<Rqا �GR��shbvk~�#x ��M��.ᬵy�����L7�oa(􆿳���2����.+w�7�@�Af8�ٕ��(�W�!Ċ&���I�JZ���+�J���q���U��@����gG���U�\ʭB��2�k1�h�H��*�I�JZ!�`�(i3�d�٣��c�A�L'��$;-,�J�d�@q�2������}°������R�wX��}�
�?�Z�,��#�2
��e�������m[�LEE�S�_�S�
ut�q���U��@����gG��y��O���{�6�*F=ॵ��@xзq8�Ј'���Xw�j�7������1H}�ɐ��/��HM���#ga(􆿳�)�~��^�~�9�>��#�DZN7�{��|� �6+^=N%����Q�K�5OoL!���}/
;$�Z��"���t})�}�
�?�u����p�����+X��FJ���-��{�"�,�>E���]�!��[@�zZ��g�f�kN�ı*�7`����\Z��K��4����/��+w�7�@�Af8�ٕ��(�W�5���^�.O¨�����+�J��Y�{'%s���gt�͓�ξ���I��RhF���k��76����,D3�.%�P;˥�'ܤ",����^�� �YW;C��K�ŶT���d�٣����Qq�M��H�_�ЩI4��欱���j���~(k��V�Ρݾ� Q2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl�ܝ�v�02+�j�V�-2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcep�y�G/Կ�]�؈9ϒ<�3$d�I�v��]huP��/��~�_Y-�<���������dC�5g����w��N�KW����rS���,�[p�M����_	�#-s����J�~AW#��WC�ڃ�P ��*����	�� ����\�'7>�W��	2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�% �t=���GR�D^;d9ךp�+�n�)D�ʵ�b��6���6�� gWVbT+踫g(�r�N�ǁ�f�TpD��ZOU;��|B����ɠ�o���3�Z��(����5���ռ�j����)w�n��ukh��MC���d��R�7h�,b0V�u�Q�ݚ�Н�A�sxW�O�Ji�];���ss2����`�|��K�z�H�MPq6.O��S�푈��^̽1��H����8�K�oe��!�`�(i3ct�:��REvє�&���ct�:��RE3z%�u�܆�#�-�p��8������aP��k�= ��j����X�u��
)\Y����4MT2g��H#�"8����{��¸�m�B��d���m l�o�1#V���<�dv��oTN֢&@��&9��?xs6'�u�&���ݠ�s�f�u_�`�ݚ�Н�K�\7}�W,�:��]]t[��m�U��Uy�~���2��}��4���,�V5VM�d�x�8�� ��ݚ�Н�$���]׽��:��]]t�L�t��n�
�s�u(�������X;p`�ϟ��7�4�.1p�Y,+
���Q�"���Urܰ#y��B7Ԅ��Y��
�iCTl�������l6��\�LtF��c����ҧ��j� �3��Nl����5	iqɍ�����~Zx�.��c�9ʼ��$ii�<�t}5�O�%E#Ps->m�9V���tpr����:4�f�Nd+l�Yҽ֗�����ڀS��d���!i�wӨj]h���6�ü��k>B2��$Jf���+��@-�-'͏������ӳ3z�]�������%kR��������֢&@��&!�`�(i3U��֜��3!�`�(i3�)ύ^��R�^Ƒ��f�?ǉ�=��){�Ysy�t��P$u��&8�,�p���ꜣ��ZLN�	��$o#[�L\!�`�(i3^P��:w0I� X�1���Õv��9e��/�7�!�`�(i3�2*Q=F�k�mD#V��A��`-!�`�(i3$��:�e�h�Ϧ^c!�6 �ef�&�2�����_�������� "5�]!�`�(i3Y��
�iCTl�������l6��/��@��:$����z�����	�;�ݚ�Н���ɕ�eY�����w6YmC,igu!�`�(i3��_(x��`�:��]]t�L�t��n�
�s�!�`�(i3p�n���:��]]t�GR�D^�6hg�}�fĉ>99��;��|B���~��D���'$c�{��lq��Hhh�f��}�� ��`n�7*�7`����\Z��K��qb	��G��W+��W�����ҧ�GR�D^ ���?R �ϟ��7�4K�ǟ
��)�;b�-�2�V��	��y��ڇ����Hhh�f�&�xW�>$�`���*1w�R���y>��yС��%G|��!� �1����p=�6��hЗ
H�ǅ��$���y�c)�h�<om���K���̂���Z��.�`��ai�}#�U���b�N��z�+�ϸ�i>hw���k$r�t�}iV��	��y#5d`2�,���l�1v] ����,�ǰ2�?~��&ĺ�����pT6cwJ��H���%�#�o����q,� L���s��$�Z;��|BljBtV`1&�\JG8:B1+D?���$���y�c)�h�<om���m��!Y����Z����1�<�l� u�<�i$D�V�"φ��<�6�@a� ��fFMqlgC>��Ӛ��S�J\7CZ�zk��Xl� u�<�10/|
�~/����l��A(�c���_G��Hb� h�ҩ�,��G��zł)w������U+��_�%]n9�K7͍��|��W&":�ݚ�Н�*qA����6\�4�@�� �-j�1tSjv�����l��=�O�-v�*_�mS8<�n�ݚ�Н�,��G��zł)w������U+��_�%]n9�ϟ��7�4�.1p�Y,v�)�DZ�ϟ��7�4�.1p�Y,Q� R��Fܑ��y���8���/�DY�7f�P:��z��l �t��D[h�ł)w�����3u{��ߤ�:C
#!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rG߸��S�Ȍ��7���9x9ջ(���'z��F����,�ǰ	M,��rER?ka׍낻��k�1v] n�,�b��,=��&(�X@�,{N�th�U�CL�ZLN�	��?ڄ��5�O�%E#P����ҧ|��sQ�G�O+�|���X���|��sQ�G�O+�|��9˫3֒�g�)�I��ł)w����ʮ��?G�+5�4��c��W������&�K�VFHN��R��?�d���&�x�����<��jkP�lX|۸Ͱ�Ǭ�j���Ÿ���φ��<�6�@a� ��fFMqlgd�G}%����3f���K��M��lak����|#HK��A(�c���_G��Hb� h�ҩί�� ff���^x��G�	B饨D���my$�N��o�/���;�Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н�y�}�6f&rG��Hb� h�ҩ�;�x'_|~�ܦ	&�P��ۥ�Y�m��6J�Ko� {�Ӻ���6J�Ko�i�Ϯܑ��y���8���/�DY�7f�P:��z��l �錛�%`��=��d혮z��l �錛�%`��c�'>���}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M��hb�����Al+�H��� ff��2�o*��g�)�I������A@�Q��ǺΕ�A�m�(�Jٯ�n
n�,�b���s����R'cf��6\�����Y~�y�����[�?�d���&����*y}e3o������(��gb#�o��_�Rv�䩲$����tb�����+�^n=\f�5>��"��qv�;-��]�Oh=!�`�(i3�'ž1�|�'����u��r��Dw\����!����#��  ����'K7͍��|��W&":�ݚ�Н�*qA����6\�4�@�� �-j�1tSjv�����l��=�O�-v�*�Va�irϟ��7�4�.1p�Y,v�)�DZ�ϟ��7�4�.1p�Y,Q� R��F-�w���+_�mS8<�n�ݚ�Н�;�x'_|~�YlԘ=��>�暩�͍΄gL;��>�a���ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ��׹����{�8�4�����V�:�RV��	��y ��f"�h-zL�EE���w����s����IX0F�MV�ҁGG`5:�����+�^n=\f�5>��"��qv�;��A�Z����r$ɓǃl[�Ƶ�1tSjv�,��G��z#�r��8ߞQ���l�N�����K����F?�{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")u��r���s�Yls��8��GMٍ���ܦ	&�P��k�Ӿ]ܦ	&�P��UB�I'���tj/�՚�-����!�`�(i3ϟ��7�4�=G���:���Y��)�D�YG�9C&��b��mf-W�c�h�5,Wlr�r%)cA �o�X�HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ� �Q$j�ލ�f���Յ.�g3ZrZ�0m�\��8�:���=���%�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��������G�&��>������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��t�o������P�����
T+Fb%��C��:O�����=�w�����5�O�%E#Py�y�Ż�"�_�0��(����5�?�J�Ń��ɖ�2i�螘c&#VL�^^J����S���� "5�]ޥ0D��/��=��K���0P��h�5,Wl�/�O'�=�J��a�U"�SƏw0�������_�H�f�M�&�;^�6#9��u��n��ݚ�Н����Y�l, 	�I��0��:|z:;�<%�a���(��	YRF!�`�(i3ct�:��REa��ZAδ��כ��p�,��L����+�t2�0�趦���o�Hc�U0�!sH�\�:ê�_���9Н@������j(2z�ܼ�P��������^��`�3J�V����U���@��������=��܄�H#�"8��!�`�(i3;���[���{s�ܱ?'�=|-�e1|E�A�2�1#V���<�dv��oTN֢&@��&���Mڷ�21!t*x�S.!ū�ez��k]m��,�۞��	�rVu,� �{k�h�+|�c�$�t�]�;���VС���u_�P�v	��YY��
�iC>N0Θ��ݚ�Н�bs��2[������	�;�ݚ�Н��Q}mҁ�t����sdb�\EX1���֠5�v{7!I���6�{�Pe�E"�I�;�q�h{b62�tstJ��:����+0$�oI�K��S&ϊ�`�y���z,3����:�v�7aaP���h���4��Q$�N�Vwk'��5�5�Hb�<�\^�
�]�xF�$3i߿�x5��vQ� ��8��;Yv^��8Ǆ1��HNԢ��e� ���� �I4��欱���j���+#c����nS�3�ǻ��d���!iV�Ո��!�|_@��0IЫ�Is��+�ϸ�i>hw���k�:5A��pw�R���y�sL]~ц��8Ǆ1����e(Sz�w��'�L���z���_ΩI4��欱���j��������my$�N��o�/���;ЈH�����E���J���U��+�Xa�H(�˕����,��&e��0�U+�qbp@�HN��R��?�d���&���W��M�[�Ʃىwͬ����B��\zF�V���P�	�#�=��R-��#U#��F:җ�S��=�w�����5�O�%E#P@?d�s�8K,Q�\C�8�Hj\��gr�d-��Z鎬�������(���=y:|}֘귈nIg�R݃��x���g��U-�e�,���6+�}�
�?�G��-�HG($R�i�Yl-�"�k� ���q���U�x��7��0��jOT�B���Q���X��+M�j�/l��I�m�d�٣��c�A�L'�O�({���p~z�r,�L;Л��*��/qRrŵ=�C8|eյ[+8��T�T�y�8�Hj\����޴��Zڥ����Ⱦ�Ɔ �����Vd��C}�� P1���~!�`�(i3!�`�(i3{�d"���ƍ2���lĸͰ�Ǭ�j�:)�
�9��W�&]�6�o8:4�I���c�90B3v�A��d�G}%����3f���K��M���i��҉)ެS��B����l��A(�c���_G��Hb� h�ҩ�;�x'_|~��Y{�<���)rl�xSNF��nF���<�W�.�P�	��
�Q�}Dw\���B���Q���X��+M�j�/l��I�m��nF���<�W�.�P�	��
�Q�}�߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3�$XR�QܛOcOZail������&G!�`�(i3�T�T�y�8�Hj\��9��T�&G��-�HG($R�i�Yl-%�z(�~�:)�
�9��3�����b�������Cҷ��e�A*�����b��Bgj��i�s�!�`�(i3��j�4�/�0���p15hQ�SQX�����RZ��P�k��!B>gl�7[�׈�m�q�/�<J|W���!B�"��ݵ�Q�n��T�\ ���H:Q ���:)�
�9f�!�Wm���m�q�/���e���W��V>�j��b�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ��׹�����A�;����v=N�]��V-[J��N0�.�`��aif��*��]�J>a`|ܘ�h��"];�.�� ���j�3�;�?�d���&�VA�ڦ�c4nǈIܺ�֝�7��ư�h-�o�dz��Ռ��W�o��ݚ�Н�b8IU_h�U���H^���R�}vJ^&�)~~;��!���c�A�L'M�M˫ɒ),��gĄ�� ���ń��	j�OpT�v��1�.0�bɩ���8�; ��8�Hj\��ň����L��b�S]O�lK��^?���+����$��r����!�`�(i3!�`�(i3!�`�(i3!�`�(i3i��r�+�<�W�.�P�	��
�Q�}FwZNE�����A@W�/�#+*f�L�t��n��}Dq�f�)�{6�U��'�U$��Y�~��k�u&����A@�|2;$�JأͽgF"?f�Nd+l�Yҽ֗�E�����+T5�O�%E#P!�`�(i3
S�z�Q�b?��t~˻�M����dN�M���I4��欱���j���MZ��;jI����aR�!�`�(i3����,�ǰ?%{B��0B�ɺ�c��5=C�Z�Ұ���,��<I��)���W�w��fD2m�O��{τ��<wȹ�k��Y@��5�Nc�X�����~X�&_ܑ�Y(�����&� &��( a⣃_B7�}�!����nސ�ш�A_�u�x�y�Zgl-�g�E�g�������(ӈ���m�r����m�ڨ�hծ8��;Yv^����j�	l@�.}�uP�V5VM�de^�~�[���>��B�K��b�S]O�lK�������[$R�i�Yl-1�*��-��4�1���~!�`�(i3!�`�(i3!�`�(i3ϟ��7�4�=G���:���Y��)�D�YG�9ž_�F��e�<Q����ON�Cf�Nd+l�Yҽ֗�Wꏄ��H���7Ә�79cKAW��R.+�T� RZ��P�k��!B>gl�7[�׈�m�q�/�<J|W���!B�"��"rH{��}TҌ5`��K7͍��|��W&":�ݚ�Н�&�z���@h$x���z(��/�h��L���2��nF���<�W�.�P�	��
�Q�}`���*1w!-㫓LT�EX+M�SU6гd��<��l�(��ԋT�W3:�h���Se���7�}�!��-��ټs�6QK���1>�n��-��u�U���(��/��z�G*�C����Uh1�;��|B���r����8��;Yv^����j�	l@v ���\{�V5VM�d��m�.j	��}Dq�f�HN��R��?�d���&�����0�9��t�P/oz�
�:qEpV��	��y$���/`�R5Q
�!`����A@ž_�F�'�U$��Y�~��k�u&����A@�|2;$�JأͽgF"?f�Nd+l�Yҽ֗���m�8lT5�O�%E#P!�`�(i3
S�z�Q�b?��t~˻�M����dN�M���I4��欱���j���MZ��;jI����aR�!�`�(i3����,�ǰ?%{B��0B�ɺ�c��5=C�Z�Ұ���,��<I��)���W�w��fD2m�O��{��JKl3y��}�	76�&�;��|Ba�&�)��H�8�:����\� ����o��=�U-���c�qDrU��*W�q_҂T�q�w���r�&U������G|M���Xr��,��d���!i"(<K�'P�2܌�B�ja�M)ikZ!+�[�x�X���+���LQ�wo��Z��Ac<�p{�5�O�%E#P��.J7h��C�x!�H��Ex4*QZ���>8
l]]y�1�b�'Be��sߍTl���g��b�I��)���W�w��fD�g�9��,Y:�{]%s"(<K�'P�2܌�h,\�NyV��FU��9T�v��1�5x|���MM
��,=?�d���&��ݚ�Н�b8IU_h��Rhy�������D����u_�*5o]Ẻ��%>�rG6j�"Hs�ĖYS⪞mf���E�i�m}66j�"Hs�l��J�&'L& �N�l_���@������,�ǰ�+9\���������������>�ܫWEFΑǜh����X "
z��_r�e~5�O�%E#P���=J����uS�#̮y�3���;_��8W�w��fD�1�C��Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h����:8ESj���b*Q}���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h��??y�8�:�����zV���z%�/��Z>L�'��D(M&��w>��Y��d���!i�T����׭�ت��+��T����oGo�Zc ��2��	\^�N���������%kR��������֢&@��&���o)�]r k�|6�8NU�:|�������J��a�U"��SEU��wj��L$?����ߐ�*U2��53�������^��n�������������Q���ËI7��-5��5Z��=��]zŎd>&�&i�H�f�M�&�����ϲ���6%�a��O���R�^Ƒ��״��/^l1�Z���=�,���9^-���2��̪
)\Y���)ύ^��z���.Mp����nZ���t��˳3[�u8�̇i�d�?�!�`�(i34�0 L?�p���@Z�_F�k-�!�`�(i3�苇��Fe#OOJd֯��
�	?�<!�`�(i3��&I���m�
��,!q�\E��0�����?Oǖqo�_����m6(\�]���f�?ǉ�=W����GS�*;q�j,���-�}s�Z�|�X[�m����!�`�(i3+�uB;y�L�6yd(��J��9ŕ�%�]�
n{h�<�o��=�U��b$�\r� 44
q_҂T�q�w���(��ԋT��D��$m*�;��|B���r������0[��Xe ��g[���K�J��]��m�'6���;8=D�P�E6�k��q��־�W+��W�OV�<��V�h�J?�߱}\��������PE�K����/�sLXNAA�����}Dq�f�����,�ǰ���������<�MP�F�}қ~Ĝ���,�ǰ����
k�=�]���v��uC�v#N�t����M~V��	��yv�ʯʗ�	�t���P����l�6��tM=br!+0�,��
������3bQ=�3�� �֤D�A��*ȑs;��|B�'�#�zا��6S����'HY-��Yk"1/р�{:��'��F�N~YMC���d��R�7h�,b0V�u�Q�ݚ�Н���M����3��~ �X;p`�f�Nd+lJ�VeSZ3&!�`�(i3Pt�d��R	}�������O9��Q��Q��O�بeD�I��k�+9=:(�I~�����h�Q7!�`�(i3*bL�(Rp~z�r,,���9^-���2��̪U��֜��3�&8�,��w�Iſ�Κes��O!�`�(i3Vx�%L��]n���@�����T�v��1���5Z���ck�7!1�Z���=������uwТ�
�+���LQ�f�?ǉ�=NM(�n��1�Z���=��m�B��dVkLs��dJ�+���LQ�f�?ǉ�=�A�����y������i�-�����m l�o�1#V���<�dv��oTN֢&@��&��|��p�S�o@�����	�;�ݚ�Н�h�'f R�苇��Fe#OOJd֯��
�	?�<�&8�,�g�Hn7�(��wӨj]h��_--���g�_�C�6%���lи{K��n٬|��VC\�2x���ЈH����@�/�MC7z���mp"�o�%�Ucf�9rVu,� �{k�h�+|�c�$�t��R����s+��6�.��6���N-Y&yo�qX� �Ĭ1�z����ْ��4F�;��%YM�	�v�3�2������"�*o�yG�f>x�:	�W+��W�1h#����5��������o��D[�h��4o�ݪ��H��q�/���˚����Z��!�`�(i3��f
t斃�B�ӗ�zjJrf����G�m���*J�X�$����q(	�fI��)���W�w��fDv���k��/9ݦ��.�g3ZE��g�Hb�t]�<Lz�B)/D��Aɶ�;Z�6j�"Hs0vZ��ҹW�`=#�e��}�Q�� �F?P�.!wG��sg嘙�^u�� 
~�F�,���XF:������X`��w{���Z���F%�X����)mSj�Txk^��]��3R��������Vo[���˚����Z��8��;Yv^���d����`"*(�D�pq3�O�̑N�$hF ���M7M�w�ToHA �I��)���W�w��fD��0[��Z���zh�QS��:Z�����nd肈��d3���2��'B>&�&i�+#c����nS�3�ǻ��d���!i-��ټs�}s�Z�|�Z�+Ěʮ����?�b8IU_h�¦�naä��E�i�m}66j�"Hs�ĖYS⪞mf��aT��3G?�d���&�zY]�埅�A���V�d��)�(Qe2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl�܎���~�k��`���7�9 �e�I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�F�I�_
S�.�)����x���	R����>�R���mK�g+�Vr���J��:�����B�����혅vº�w�⽒���M����A�m�(�#W�U��ظ�d���!iR����
w���������q�©�����<�������~s���^��ӳ3z�]���ϸ��#|S������3[�u8�S��Ǵ��BR�^Ƒ�ӡP�Kf����|�F����A�+�~@�\��qZo����!�`�(i3ct�:��REvє�&����d�uY�ؤ��E��!�`�(i3Ĉ���rl�خd���!sH�\!�`�(i3C��[�����p��@LC��[���ԗ��6%�a������[��C���������a����"�$!�`�(i3���ȍry��	-�E��%�~�X����Z鎬�������(���ۯ���@Z�2[QvA�N��L+@���w�K�R he��as�C�G���-�p'�"�hPW���[f=HJ��nt+hjjp��2[QvA�(%�(�Y+�(���B��U��0S���NB�D�u.?;�^H���"X��[O+oF��!�`�(i3^�9.�JQ�0��"��S8�ؘ�Q�t�+�g�>U�CC����/�F(�@vW4��`�|���eC�����jA��L��)��$3˓8���/�R݁��!�G�+�g�>Ub����{����ITf��J�� m�Õz������\�����wUm�y����}D���ݚ�Н�[�л���7ۤ�ǲt'�<	: ��YC��?�!�`�(i3$���]׽�#XEXj�.h�J?�߱}f�Nd+l�Yҽ֗��"X����ݚ�Н��9+�����Rz(��g��NEP�B�iY�;���!�`�(i3k/�z�xEQ���*[UxG!�`�(i3�|�)՜�4�a�/!O�+�_0c ۜ���,�ǰ&k�����dƉ��u�Z��E��3?�d���&�F�I�_
S�0v�6���!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcۖh��)�ԯ��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h:���I�8�:�����zV���z%�/��Z>L�'��D(M&��w>��Y��d���!i\o�LCd藀�)�_f����/�sLgwe�ŉm�m�jp=�>��o�
�v}�D�~��*�7`����\Z��K��~�]D�o"ly]/�qF���ӯIJ ��`y�����n4s1�	u�ɐ���hu*_�+��T�����h�6ؖ�(����C�-�nC/$PM�^-q�x�l��1:�N�*�x���N�#,�	X���CIaZ�x&_FA"���,�7�%�a�A�m�(�S�gd���zg��p��I7��-5�B�wj$g-��W����vcyj;��q,G����?���_�\G��4�	B45Ji�];����z~~�Y_" �g8Yw��u��n��ݚ�Н��z~~�Y_"R�W�u�B�wj$g����d]���g�P�e�9�y�3�A�e����kn4@Q�/�!�`�(i3���ꀍ!�`�(i3�˺�Q���f�?ǉ�=�M�g����!�`�(i3H��bf�?ǉ�=�|�)՜�4!�`�(i3�a�/!O�f�?ǉ�=��TBd��pS�*;q�u��&�o��n<���AV2�?�+�p!�wӨj]h��
����ŗ&8�,��ĦsW�0��Ϝ��*@&+�_0c �bYގEV�tպ� ��q_҂T�q���e�u�V/=T��?�N�����H+����f>x�:	�W+��W���̈́��3R&�5�V��X9���d�uY���d5z�R��T�\ ��;��|B���r������Uz������/�sL��t`x;��wiV7Q�h�J?�߱}�'��$zөfĉ>99��;��|Bɖ!v��wm������w�R���y���,!��:ԫL�S��7�g]�[ŽV��	��y��j�}�-�	�t���P����l�6�� ��Z+0�,��
������3bQ=�3�� �֤D�A��*ȑs;��|B/B�Â���2�εp�K�Q��O�بeD�I�F���������Z�ש���&��W�{C�A�n<���AV2��O}�c���*A�Y�{'%s�[�&B�踫g(�r�2������"�*o�yG[�����ݪ��°������R�wX��C>��ӚH�RtV�^�y2Z��ZkB�@o��[ea�8����:%��Z��vDY�όW#VL�^^JR�7h�,b0V�u�Q�ݚ�Н��������r�E�Y������i��tt"���O6/��������рӚx�f�?ǉ�=�]V�H7'�R�^Ƒ��!�`�(i3 tZ�u���ߘ�)�Ij;��q,!�`�(i3�z~~�Y_" �g8YwU��֜��3����d]���GF��a�1�Z���=�,���9^-�S�_�p���it	�T�=��?�AQ�0GȨ��_�\G�k�y'��af׍�Z���e����kn4@Q�/�!�`�(i3̇i�d�?�!�`�(i34�0 L?�p���@Z��hy��Q�#<4^�-����b=�!�`�(i3�չ�Ad�!�`�(i3z�Gb��P�!�`�(i3��TBd��pS�*;q�u��&�o��n<���AV2��O}�cD�����m�wӨj]h��
����ŗ&8�,��ĦsW�0��Ϝ��*@&+�_0c �X� �Ĭ1�<^��0�u"��D5�|أͽgF"?�Q��ǺΕR'),��`�C,;�m�~�?�d���&��ݚ�Н�ۆٗ��NJ`@���!���ƫ�P�A���8��''6���;8=D�P�E6�k��q��־�W+��W�.5o�fa��N����Qѕ&D�a�Y��m�'�¯ԙEI�s+��6�.|th1�$�g�ݚ�Н�w�R���ykb>���p׮Miz���;b�-�2�V��	��yG��Γf��Bp����ӛ�i��.}�	76�&�;��|B}2_R��'3x)'�V�*�?��O���2�"��H�ʱˡ�ۿ��j����H�V�7�}�!�����*�t��v+�/;$�������1�1F%јI$r�t�}iV��	��y�bB�.�����	7?�����,�ǰ�QCT�"�Ʃ�A���vA#&��Q2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�:1j�=�+���u&Z�=��O}��� 3[Hn��Xa�����`��O��m�]wew1"G�6L_i��Y8:0nQ�rV����X8(�K&'3����G��-^/s�B`@���Uc�`X�,4�?n�J�����W���h,3
V�R���S�sq��u�����|S����	��rc����	:�¿D�?��	`��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�{zY����b�8�dX�↨q�©����y,�m��M�5��MC���d������S���� "5�]W���`moF˯�+)��h�\ƙk����p�><��d5�:�w�+���LQ�f�?ǉ�=h�5,Wlr�r%)cA7]��l5TI!�`�(i3+�'T��H����8���)�Um��T����M��6i����v(�ÂfC` ��\��u��n�:�'&�
x#2���p5�}�]���8!�w� �O�z����7�]�hk��,�:�N�*�x��0�&�ͭ�&8�,������	�;��=����t�7��r�=Tl�������l6��ƿ�d����X;p`��Ĭt�'���g�4�������YL������Y;�չ���1_�I<�N��[�л���7�&8�,��ĦsW�0��Ϝ��*@&f�?ǉ�=\.�l����k��r�a�^��D��
��Q�# 2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�$�/T�!J�`���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�Y�o��}�����k��h`�H�MPq6.�yܤ�܎~�J���^W�������������_�ft�m-���L%�o5j
�^q�&Ѣ�� ��&6�%�@��n{�\�<:���\���D)�g�%v�=̽�0Բ�ȁ��;�<�h�kIp�#J,i�~X�Z�o�x��o��ײ]�4�Kq%��M�Vr���J��:����;�	��o�g��}>�IM8e�׸J�q��G��m��+�Ƽ(��h\^�N���������%kR��������֢&@��&2�w��~)@���k�֭AQ�0G�C�`�/�t���E�����u*_1�Z���=��m�B��dIR*�fN��iGR��o\j�g��$Piq�VD�Lg�����X���ݚ�Н����8�8e[m��������iq�
�Bk�i�E?�xu�1#V���<�dv��oTN֢&@��&�_F�k-��苇��Fe#OOJd֯��|��p��PIQ#�C,0�?��ʉ��%>�rG��M���ʩG`B� f�?ǉ�= �@��&}� ����'_�D�8 !�`�(i3@ E������n�T�����+_AdVw�R���yh��7�S+���
e�l7o�V������.#f{}#k���4&Ƒ:2�c<�^<�H�W+��W�|]η���7�,��n6�o8:4�I���c�90B3v�A����èV\���F�`yx�>�+X�M?��y�!�`�(i3+�uB;y��'DV���b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3L�)9�/��22�ݚ�-����!�`�(i3+�uB;y�ڇ������ � �"!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j7&�u��F
*��q�)�`Vo����6j�"Hs?�L��4�Y]؜�t2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��OC�0����t��[���P��EC�`�/�t�KV*�3?�|��T�5�d�,W�He�!� U����z~/�}��j,NJ��:����8���SY�N�o��C�0�_E,�8�o��_�Rv�䩲$��GQЌJ
�յ[+8����"sS<�0�zG�������&G�wӨj]h�(%����K7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩ�-��)'�E��ȷ��#o�]�ʄǾH/�d��_�mS8<�n�ݚ�Н���4�*BqC��~�;ϔW򻐗�NGq���ÌZ>u�,R�� h�ҩ��wӨj]h�(%����+�uB;y���O�	���lC��U�T�\ ���:5A��pfĉ>99��A0ok�ª���l��������t�|ݔ�3�5�}�]�����nv��~���$r@H�RtV�^;�jmT�#��|�!�[�w/	��^#��4,�Q��+�uB;y6R��*Q�z�ׯ�1p1�Z���=��,�����!���2�(+�uB;y���O�	������v�h��4y��ij��X� 2!�`�(i3>_�Bnˌw/	��^#��4,�Q��+�uB;y6R��*Q�z�ׯ�1p1�Z���=�1�(�yj�!���2�(+�uB;y���O�	������v�h���ў�L��-����!�`�(i3q�\E��0����G�t���m�� �ݪ���CyW�f�tR�wX��!�`�(i3�	��x��ݚ�Н�����l��q�P�oV4ʐ�}	�[���&�ŁHL�U���W�����&G!�`�(i3�wӨj]h�(%����Z鎬�������(���/%Z�ڄ^1�B/���q%U����z~(����(]�U����z~)���	6�!�`�(i3�Ra])n#���r����!�`�(i3�� ߌ��̷_��yC��S8�>c��6/{v=~P0:Q+�3yK������v�h!M�T�ĥ��P�7� �:5A��p!�`�(i3���F��O��ݚ�Н�fĉ>99��A0ok��
�:qEp�;�P�t�5
�:qEp�;�P�t�5fĉ>99��A0ok�׹�3��܌o��oŵE=�[�P�X;�Z��;_��8W�w��fD[�P�X;�Z<0)��TG䟳��LQ�%�+2��k��kK�I�Q4p�/Cj���C�1A%^�Q��U����z~/�}��j,NJ��:����8���SY�N�d�}����U��)���Y;e�iK!���d.O.C��|#HK��A(�c���_G��Hb� h�ҩ�{k�h�+E�g�������(ӈ���m�r����̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l���{$����^V���!ֿ*Y��b"���LQ�/81tSjv��wӨj]h�(%����Z鎬�������(���[���-���W�6?��jsrCm�k#��2�bD�=�^݊��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M����m#p��ܸ2߆X�.�g3Z��S~��L�ѧz~�u2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!QY_׬�af��pD��X{�:{�f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc[�IC�r`~@JFa�i#¯��TG6�o8:4�I���c�90��G��6�(&�L��'ž1�|�'����u��r�幆i��}��_�/}	�dN�<@Iv��nt=:��:5A��p�T�n��a�M7�a*���,\�����k%�B��;���N^�|`#�BO��he�����'1�m+�D8*qA����6\�4�@�� �-j�1tSjv��
�t��T&���LQ�/81tSjv��H�����d�@���G�Y[�	���ġ��,/�r�]/2�ݚ�Н����8�2����o�W��g��Ȋ�>��������w�w:�!�`�(i3��i��}�a�E�Rq���my$�N��o�/���;
�:qEp�;�P�t�5����l��MmN}4��vI�o��v��ONH!�`�(i3��i��}��?@k�(м�{!0g|p8��"�n&>��������w�w:�!�`�(i3��i��}��?@k�(�97��EN�h�h�u+��.ᬵy���ܝi���d�@���G/��S���.F|�r����%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��j �_�ȇL�X Hz��0�Jw��3��o�c,�̄���{�=0|yY:��{�o��_�Rv�䩲$��8��I��.��|ȃ�A(�c���_G��Hb� h�ҩΤ����3�_�/}	�dN�<@Iv��nt=:��:5A��p�����3�r^Fn�$|dN�<@Iv��nt=:��:5A��p�����3�?@k�(�dN�<@Iv��nt=:��:5A��p�����3�K�?\B�]E�g�������(ӈ���m�r����*qA����6\�4�@�� �-j�1tSjv��
�t��T&���LQ�/81tSjv���!=.�
���5ʦ���*�·O�f��1.X����l���oi���:�9�qw*{c�i7��c"?�Á�ݚ�Н��)E�Y�ȕ��U�._�nQ�rV��q�t7�B� �b��!�`�(i3�D���s��l�
@\��L�溥����v�8:?�'����-����!�`�(i3Us��K���fx�	��j �oi���:6 y2��R�՝� s�#���k$ ����l���oi���:E�g�������(ӈ���m�r����
�:qEp�;�P�t�5
�:qEp�;�P�t�5����l��!��3ٯ[�8Y�^V߶�9��\��E�H�RtV�^�Jo���j�oi���:|б��4����-����!�`�(i3Us��K���8Y�^V߶�<;�ò1���G��t| ��a!�`�(i31���~!�`�(i3�����3�?@k�(�97��EN�0�2l?e���yN��7��aq��8�1��e��],��%s��^�y��� �s��c�!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�o�u����Y�$�Q��b{|�|ʫ��ď<�+��9���2�"�G�p�P�(��Iw?�d���&��*#�m z�wi��r���:�Nz�]'\gWg��	�Z�kfc?�#	*]]�(&�L�xjzӝ���I(͂��-�����'��o�/s�1��pE�g�������(ӈ���m�r�����ߎ ��E�VTҝD!u��nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h��-����;�jmT�#�,l����M?��y�!�`�(i3	�)��&ghRV��R�4br����}Dq�f��Zj���
],��%s��ԏ ���ԭ�m��3��p���H���6Sa쎑t2�������50f
V��.ᬵy���Ÿ�`u�1tSjv�!�`�(i3�I��� g�����Օ��qvdЧ^{�jMdGN���!�`�(i3�'��o��̟�1�C�|J3J����#�=3!�`�(i3�����!�`�(i3�ߎ ��E���Bf����{_8�Y��=�}�Vݨ��}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j��Zav����U�3N����JV��	��y ��f"��4br���fQ�J��� hew<�+��9���2�"�G�p�Pڹ��/^�w?�d���&��Z�֓Ei��Bf���������I����,�ǰTm�v��G��4br��i��^�t2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl�ܴ����-VL�����[�R���'+_��'5��F=<��p*e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc,���H�z�+5�4��c���Ÿ���φ��<�6�@a� ��fFMqlg{y����i�q,?5q%�d%p���T��Û�r$ɓǃl[�Ƶ�1tSjv�9�{�Jj3Ř�z��l 	B饨D���my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�B� �b���H�����Yu�������&G����l��̻�>a�8E��XE��� �GR��shbvk~�#x��q��ZVT�x�"��XƤ5_�J�	�LÆ���#��p��;�{��!�`�(i3P���x�NS���U-�y��j�ł)w���`�b?�ݚ�Н���jVѭ@!�`�(i3ϟ��7�4ÿ����Ԃ�nF���<�W�.�P�	��
�Q�}HN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}�~(����ϟ��7�4�Zcd��Ԗ�ۄI��K��p12����2{i�����s�;�9�����:�.�赒�-� a⣃_B��!��8��&��@ �'���ȇφ��<�6�@a� ��fFMqlgd�G}%����3f~(�������u`�`J�A��xjzӝ���I(͂��-����.�`��airV���qޤ%�n#� �nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h��-����;�jmT�#�,l����M?��y�!�`�(i3P���x�NS���U��í����+5�4��c��W�����+���*#nC��6�g��z���7�a(􆿳���ʽ���~rV���qޤܡ��F؝=��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�MR����}������+��;_��8W�w��fD���u`�`�Zcd��Ԗ�u���bΤ�tA�Ɏ�A��朢֛�l����c�n�RW�A�&hH\+��O�r!�J��:�����V5VM�dC��6�g��x����K�my$�N��V5VM�dC��6�g��``�^��c����,�ǰTm�v��G��u`�`�Zcd��Ԗ�j��A�ؼ
��ь:�Gɩ��IX0F�MV�ҁGG%4vkz����`���φ��<�6�A$�ʁ� �o����*�'ž1�|�'����u��r��T��{B�z���b�z)iŞ�W�%3AԢ�a\�Zx�.����#��o�TX5Ȭ7�j�W����^��D�Ϝ�}Dq�f��ؼ
���O�k�����nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r��܌;���'����u��r�妷��ҧG9�:Q��
ϛ�(L�p8@)y@d��{��1BWW/S��8(�E���Kt����ӯIJ ��`y����ݚ�Н�;d��'�XƤ5_���H(�T�O��{Tɀ�"'��&އ�[t�Y81�d�@���G�X���.��ġ��,l5R?}�b����n)5,�O�޳!?�R��n}�����H��B� �b��!�`�(i3#�+���?}G9�:Q���'"�8�5�� h�ҩ�V�Ո��p8@)y@d�`����n���P�|TDqId�ja�<om��h�a�'�ȷ�H���9�ªe`���1�m+�D8
�:qEp'{w#/ B!�`�(i3�ؼ
���'\��i�`)[�-hnFX�``�>������fĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹���C���N���]J�oW��`{�n5��=�ɟw��D�����˦G�G���۵z p8@)y@d#�أ��+����,���N�����x��t"�ؼ
���$����G�ش�oh��a?H9�v-Q�WdM4@Ȁ��0��_Թ�,N��1����l�ˮ�N��j2�K����S�p�d.t@S�MgW�6�h�g�t��-��4�1���~!�`�(i3!�`�(i3"(<K�'P��ƣy
���b�Bϱ�nQ�rV~ù,�u����7���{r����������X��3�BS}PR�]C$�Jw��3��<*���h�>F۝��k]m��#���6���2�"�G�p�Pڹ��/^�w?�d���&�Ms�����x��c�ۡ��W���\��'���Xw�j�7���ؼ
�����b]����m)�X�\
ihc�ؓ;)05 S�s�lZ鎬�������(���Κ^�q 
�v1a{J�M�ld�zPk��!a�tc�&ck��°������JB8�^C
���;_��8W�w��fD3 �����}c��ko#��C�eݹ�,���H�z��ݠ�s�5�A�)��?��u�h�5,Wlr�r%)cA��z>9�R��d���!i�[ie->fN�2[QvA�r)1;�Os�rs�i�E�8�w������5ʦ���.J���0z�cULj� 1�B��/����9-��g���t�
�:�WdM4@�r)1;�Os�rs�i�E�8�w��ӗ�"��I\��! c�A�L'4��"�����WdM4@��hd=��&q^�`
�c��><�$��;mQ��8���/���/z*x�n;��|BE��Vˀ��e�8�ʫ�ޚ��Jt����J��4�5��tA�Ɏ%�<'L�+��T�����D3��\^�N�����ϸ��#|S������3[�u8�U��֜��3!�`�(i3�:��]]t}c��ko#����z��,Wc��IrM�e<�!�`�(i36�X��U�o̥�0�L�p~z�r,,���9^-�ss2����
)\Y�����'u���ɿJ�ҧ{�x����y�mZH֫&��5�q	�gh�䊉�䞘gx�n�W�����v;�k�@d���t��˳3[�u8�k/�z�xEQ���*[UxG�y��j��k
e�3+{�i�m�T�੉��%>�rG��M����{����"q�\E��0��n���Î��ݠ�s�M6E]s��?V��j�c�;J�*%nߙ���"���t��4�"���S�;��g-�:�Gɩ��I�?g�f&:��r-,N�[8j�cR�7h�,b0V�u�Q��M�=�@���k��!�`�(i3�N̮�$�WdM4@�_B��f�?ǉ�=�gCu(o?C!�`�(i3y�Z�;���>0�1ۍ�h �=�f�?ǉ�=^P��:w0I� X�1�;LV^Š�r��Lo�_jo���po�h0�h�#"
s���
|�1�0j�$��:�e�h�Ϧ^c!�6 �ef��BA�IH���O,8��=����t�F�,�U6�Q�L��֭�h��O5�tx\s�l.�	�C���ɕ�eY�����w6YmC,igu[�л���7��+���ihc�ؓ;)�<Z�-q�\E��0�]��8ƹ��y�H���7�el\wG�~�פ2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl�ܴ����-VL���������P���d�Mq�F=<��p*e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcr�r+�� �s���〼� n`Ip�`,9�H�W��`�z����k!�M�Z���	qb	��G��W+��W��Ɔ �����Vd���ة�蝌b�Bϱ��Ɔ ���	�ϝ�YC���;_��8W�w��fD�Ɔ ���ڣ��>7�s���MS�:�GI�^��T`/���혅vº�w�⽒�J�	�LÆ���#�喩��H�V�n8�A�A�/�����sc�̆�!Y2dyӣܡ'iŞ�W�%3AԢ�a\�!;���}�ߜ�*�l8�b(�����-\71v�<om��-T�"�N�i;��#��F�r�f�tm�;���W����G�iA'R�	��ೈ}�β3��(6]���P�|T|o��M<!�0�=<MW�-}�	mpTUÙ���#���FZ!��9z����9�9:�{q�����i���A���;_��8W�w��fD�Ɔ ����x�-.f��F�J���ى�zա~��M��D߫�ܢ	Ϧ�s��,��T%���a_�}��0ͅ�f0�	>c ���l�I(/2]�;�6*���z�Y�]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7r��*�tZ?Zaze�oY��˿^�S�>�������"sS<�0�zG�������&GЈH�����b�'Beͧ��&�~L��8ƿsE�g�������(ӈ���m�r�����nސ�ѽv1a{J���ǔ���'�P$��!���?t��my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�B� �b���H�����Yu�������&G�B�'��a�/�����sc�̆�!Ym��q,�D�z|5��z�C�x!�H���J��Ӊ�T���j�7��}D8_)'!��r��ݚ�Н�N��	�Ȓ{A�dha#4\�0l���8ƿs��DKY���k]m��F���d H����S:Xң�dC�m��3om��:5A��p���F��O�}�	76�&�� Ӗ�t$�)�vx�YL�P��tõ���lF���d Hm�q�^�g�Ɔ ����;ƹ��:i��DKY���k]m��F���d H��(әaZ��h���S>4�mD �d/Yڧ�;^�6#9>���@]"X;�3/���k]m��?�Bo����Ɔ �����O�����C�1�r5��(әaZ��h���S>4�mDK�?\B�]i;��#��F�r�f�t��s�P|~-�;ʾ���j3YY<r�!��'HY-��
�C��n�%GV��o5]�Q;�im��ȍry��	�
�I�>y!�`�(i3��i�\�{q����W�Ty��5��){�Ysy�t��P$u��&8�,�oa�}��p�-�o%�݃��x���Ԓ��t�2~?�������g�����t��:ҹ���7��I������-5Ԥ0Qo�n<�!s
9��
ss2����
)\Y�����'u���ɿJ�ҧ{�x����y�mZH֫&��5�q	�gh�䊉�䞘gx�n�W�����v;�k�@d���t��˳3[�u8�k/�z�xEQ���*[UxG�y��j��k
e�3+{�i�m�T�੉��%>�rG��M����{����"q�\E��0D������'���Xw�j�7���Ɔ ���9/�^Â?V��j�c�;J�*%n��Ɔ ���	�ϝ�YC�����%�!���Gg�&�B�~�aV~����E�+��@-�-'͏���������=���t�iZ]XF�hx��G�����Fz�U��֜��3!�`�(i3�kޮ��n���㬺����<�����"BqYr�X�<\�!�`�(i3�����
L�c�n�R�HM���#gmB�z�$�~?�������g�����t��:ҹ���7��I������-5Ԥ0Qo�n<�!��t&�"��ΡKCh��(	�G��^����K�7����&Y��V�s�p�˲=$��:�e�hfH'��!�i����VZD8X�˞�DG�O�G?X2�K��2WI'�=��y)k��>���t��˳�O�����M�g����H��b8X�˞�DĠi�d�?�4�0 L?�V��=�4�6[��u�9k�\,���a���&s�q�\E��0D������'���Xw�j�7���Ɔ ���.�&�?�����X��{k�h�+:A=�O���C�x!�H����0pJ\�<��E���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�������'�al��p;��|B/�~��,�����~�k��`���7Ք�)�"e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��CNK��v�n�2)F�eCo����q,� L���>�"�x�׏��Z������23��
�
��(3�� L+��"��ӌ�r3 �����|���|��B�R���$]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7N2��j������mA�7�癆cgQw�c4~Nr_�mS8<�n���*y}e��VU[���I�)�ݳ���b+}y[�k��^�1��dc�@c�����h��-�����s�Yls��8��GM��-����.�`��ai��NEP�B�ۥ�Y�m)���A7��!=BM��~_"I�����.�`��ai��NEP�B�΅i�����T�B�X
Ŋ�0����g��U-�e�ott�i ���NEP�B�΅i�����T�B�X
Ŋ�0�����"X��[��I/J!�`�(i3)���A7�a�@����Àg�)�I���T�B�X
��j��8�u��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6��������T�B�X
�F�Q�f�)IA����Cj����tL(�g��$KB[DA���hvl��9�h �=������-�S�h �=�*�a"4̥�0�L�p~z�r,��:fۇ�0�=<MW�-}�	mp,��_А#�<om���Ϻ� ��H����8�(����������cɧ �GR��shbvk~�#x ��M��.ᬵy��	ۢ�wz[k��q��־�W+��W�fePh����X2UbP�I���x�a[M��1�:�Ω�����|"��YO�.Ŝϸ��#|S������3[�u8�����$G⃍�������������;^�6#9��u��n��ݚ�Н�rM�e<�!�`�(i32�ln�_It��9j.�l>'�o��&L�/<�t��Cn��P)��	�+�`g�]@n_���?3".3�]�N�L�溥����v�8:ۛ@W:���#���F��*{�욋�Օ��qvdЧ^{�j)�]�T��z�**ߜ�*�l8�b(������l__��E� )�&��,�~ ���@1z�+J���5���Adu�5k
��Fɴ|�O�j�gh�䊉��	��J�6p�N��2��,Wc��I$��:�e�h�Ϧ^c!�6 �ef�&�2�������ȍry��	Y��
�iCTl�������l6���0�&�ͭ�U젩`#�4>?� �1��ɕ�eY�����w6YmC,igu?V��j�c�
���!8Z鎬�������(���'�jh�,o�����S!�`�(i3@ E����8c�j�;��O�"�\� o~֊&w�R���y�E�6������=b��uǓk`���)���1�J2�*���fePh���� e���K�_�t ]�,�����}>p~z�r,؛��ap~z�r,k�@�&��T:5�����2������}
���!ꭶ��yN��7��aq��G�n���t�;���NI	��y7DT?�R��n}�����Hو����w/,�L�溥����v�8:ۛ@W:���#���F��c��k��q��־�W+��W�fePh���� 2�:����]�!��	Ǹ�y85��J����;#b��?���;_��8W�w��fD�{<_�S^��Z{oBQ��;��O�"�
9�S�F@�����jֈ�U�d�#�b��i0c�������D�_�k�W�A�&hH\#j~X�6W�A�&hH\���2*CA>0�1ۍ�h �=�Y�Eb�3��;�WQ�.p�2������}u��Kh���m��3��p���H������7Pr��ġ��,ˌ�����'�̗����Qnջ�%�f4�����p���yN��7��aq��G�n���t�;���N�b=�)3 a⣃_B�h���Q�kUx���6_����kY�O�Z�_�m��+�Z����y�MC���d��R�7h�,b0V�u�Q�ݚ�Н��
�I�>y!�`�(i3��i�\�{q����W�Ty��5!�`�(i3�gCu(o?C!�`�(i3LZR���[������2������}F�G���d2������}��s�5e��g��cH�wA�?�p�p�{V'��kd.Cf����+9��lE딧 �GR��shbvk~�#x ��M��.ᬵy��ݼ?����DY~�y����o)�T*�c��n�da�ۣ���(�犽{Tɀ�$����nQ�rV,?�����k��M���'abW�5�}�]��ϵ��t�pu:�]f�?ǉ�=�O�G?X2���Y �6�ZWq�ߑ|�ݚ�Н��W�"�Ů7�6��,�ݜt���,\ͨ܉p����O,8�ݚ�Н�h�'f R>N0Θ��ݚ�Н�Gظ0����t�%�Z?��<�ry^�%��C����\P�ʊQ:��IK��<[�л���7M+э4��Y�{'%s��jb�ܳ�/�����b>I�Wkxf�?ǉ�=D�wP�/�w���bc��U�d�#�by��W��;_��8W�w��fD)IA����Cj����tLB�'�4V�������� �a���GE���T��>f�l0 ��J��9j.�l>'�o��&L�/<�t��Cn��P)��	�+�`g�]@n_���?3+��y(��'{}yw~�귈nIg�R�5��/dV�L�溥����v�8:ۛ@W:���#���F��*{�욋�Օ��qvdЧ^{�j)�]�T��z�**ߜ�*�l8�b(������l__��E� )�&,�W�8"M�5�O�%E#Pڗ����7���T��>̷_��yC��S8�vV�y��F�k]m�������%�w�R���y �+�5�?+�T��ˬ8��� �r-��M�s�����%8&�d�I�_#�	�Zz/3>��-��k�5��05N)hiW�U����҉�p��P���x�a[M��1�:�Ω�����|"��YO�.�t�iZ]XF�hx��G��N����p$��<
DN͗&8�,�nU�gF�r�f�t���MK�L��.��֞�������i�����+��c_�B&��p�)Y����2�Yd������.Cf����)Y����2��L�溥����v�8:��|`��'J�	�LÆ�c�9ʼ��$�G�nJ `G�p�P�F�����1�׀���ץg_�,���+^+�CǘHs��BQ�~k����C�x!�H���f񓟗������;�1kT�|o춍���m�s
9��
Qov�䆙��K�5OoL�H��>�9��'abW�5�}�]��ϵ��t�pu:�]f�?ǉ�=�2*Q=F�k�mD#V��A��`-�K�^����\_9ͫ��Q������(���^����ȍry��	h�'f R>N0Θ�(�6k�4d:$����z�����	�;�;b�-�2���:��Zg�Hn7�(�?V��j�c�
���!8Z鎬�������(���'�jh�,o�����S�2��}���zgm##����Н�����r�s�����%8&�d�I�_#�	�Zz/3>��-��k�5��05N)hiW�U����҉�p��P���Q)�+J!�1�:�Ω�����|"��YO�.�t�iZ]XF�hx��G��N����p$��<
DN͗&8�,�nU�gF�r�f�t���MK�L��.��֞�������i�2���|Q�c�n쯎+�ܼ�P�����2@�n��j(2z�ܼ�P���#�紩$�_�B&��p�)Y����2݃��(�犽{Tɀ���S�<Ԣ�E,�J�|R�ZLN�	��D9������G�p�P�F������c;xć�&Y`��!�z�-���1��C�q��A�c�b�'Be�m��j�5�d���I� ������B�>w:] q��j�J^2�Z���8f:ҹ���7�`
�����Wss2����
)\Y�����'u���ɿJ�ҧ{�x����y�mZH֫&��5�q	�gh�䊉�䞘gx�n�W�����v;�k�@d���t��˳3[�u8�k/�z�xEQ���*[UxG�y��j��k
e�3+{�i�m�T�੉��%>�rG��M����{����"q�\E��0D������'���Xw�j�7���Ɔ ���.�&�?��B7Ԅ��p�n��N�Sm�@�<_3GH�F����u�ķ�s+�d++~l!�$�"���+!�/}�`,9�H�W��`�z��Y��),�B۸����H�V���!��8�䱬s�^��\�y��d���V|���أͽgF"?���(�犽{Tɀ���S�<Ԣ�E,�J�|R�ZLN�	��]�F��K�F�!��c�N
������Y�U���f�6l�}���)d�F}���V6��b�g�~.@-����5��] 9�s��M�ߜ�*�l8�b(��E,�J�|R�ZLN�	���}��~_�w�;T�^W���}���i���!_���'F��&d,4��6	����ҤyM�d�X�\m+)�15���P�|T��D�?��/��j����?zk�8g��mT�Of���-A�¤�x.�Knq��H�����ġ��,a��bt��#-��[�xw=�K�G��&1���$�yp|�,���yN��7��aq��͹��e�[�.ᬵy����{!�)X+J��a��PƐ����r��������]�Y�_�H����z9�9���K��T8��4��L�O]'\gWg��	�Z�kfc&�2������èV;�jmT�#bs��2[�a��o���H�RtV�^��k�C�-�<�ao����O����8Q������51�X�c�rs�i�}�O��L��_
�uk*����S�~���e�)qP@L0��U���(�犽{Tɀ�$����J�	�LÆ��S1�c������b5?H" 1����>E�%��*d��:=�;�մN���_�Gt�7A�;�֋`NY~�y����u{ᵿ����ݚ�Н�=3}��~;=��X��/�-oRCGtKż����51�X�c�rs�i�}�O��L��_
�uk*����S�~���e�)qP@L0��U���(�犽{Tɀ�$����J�	�LÆ��S1�c������b5V��$@C��y	����F��،M�Rh�O������ڽ��^̽1��H����8��ӯK���
�:qEpk+Q�h'�Ȝx�5W ��̫(� h�ҩ��H�����Yu���*Y��b"Wfי�b��}!D̅��}���wWfי�b��}!D̅����A���HL�U���W�����&G!�`�(i3x�&Hg 35+�L�^� h�ҩβ��y��lDR�6؄���c�ۡ��F</h,��.�W	/g��6��c�ۡ��F</h,��#m�ڧ[�:5A��p���y��lD{<�)��!�`�(i3!=��+�Hb�2�Ǐ��Pn<����I��i�h�]�� qY�{'%s��n��(��n�v�ĺ�֦�w�#d�y�=�����!�`�(i3E�xa�/ݺ�A0ok��!�`�(i3��KZP2D^�uPϿ.����"d����Ľ���=B��7��i;��#��F�r�f�t#hԇ�H�RtV�^!�`�(i3,�0��J�������+��<�ao����O����8Q�����h��g֕����/�Z�k�ʆ-�(i�pY%���m��3��p���H����HRCJ��<om���o�p��F�����+!7Ev-}r��C�r�X8g��mT�Of���-A�¤�x.�Knq��H�����ġ��,a��bt^��9^�����-/a8!�`�(i3�q�9�ͭhy�`�w��v1a{J��\>Pq�������B]�PZ鎬�������(����.��$�ʸ%�])�+�}c��ko#��J��ӉA���m��i���#7X=!�`�(i3�Ra])n#���r����!�`�(i3I&!y'}�}c��ko#��J��Ӊ��K��i��̷_��yC��S8�͍u�	�g؝�b�Bϱ�]h�(NAP/i�\	t�R��-�g� �GR��shbvk~�#x�l7�l�r�#���F��|}�&��3���.1t΀�+I@Lv�@[�JJ1��P�M����jN1]�U����ڽ��^̽1��H����8��ӯK���!�`�(i3fĉ>99��A0ok��!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ��׹�=� @������1�sB:�cV��	��y ��f"�I$T�w����	Wa=�h�i>�Oi�-4m�TF-���?4���R;���t�T��?E-h��`f���sC>��Ӛ��S�J\7�@�f�smy
�߲yR56�S��M��rs��xjzӝ���I(͂��-�������%>�rGWfי�b����{�6�9\�B^6�/.�<����㾸b+}y[���%>�rGWfי�b����{�6�o� c �"j㎡(�%��v��!�`�(i3v�A�
^^3�V�C��k�&�c���f�s栿o��$�\%e��}Dq�f��L�����B��2�k1�h�H��*��s��Rm��u/�Ο/��kOT7�wtMM�0�5G,��Gc#i%r^�����8<�l^�%��v��!�`�(i3R��ak����`T�ҩ�	r^W	��s��G�z��%��v��!�`�(i3R��ak����`T1�h�H��*������A��b+}y[�߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3e<�Ia��la��o���H�RtV�^�6[��u����@~H�k����`T^X�eg;�5�[՚1DNh���W<˥�'ܤ",,�����;	Nh���W<˥�'ܤ",��o5�����,�����!�`�(i3��9��稕/Tu���Ŝ��%ٿ�ˉB��5��*@����Nh���W<˥�'ܤ",��E� ��"U�7s,�/Tu�����_&������@���P�d����%>�rGWfי�b����{�6�o� c ��~�����U�s
ƺQ׆��p0�Ĝ(�IyIR�%r?�	rWfי�b��}!D̅��t/)������&�K�VF!�`�(i3�L�����B��2�k1�h�H��*��s��Rm��u/�Οq���3��`��R�`��ƍ � w�u"��B��2�k1�h�H��*x���0�
&YY��!�`�(i3g�>x�����H��6��b�4ƭ,�t��2� �צ�L��^�뢗�˯��Wނo̒.�9�lA�J�����7�wtMM�0�5G,��Gc#i%r^�����8<�l^ܲ�}�%DܭD��_�W�.��;�#�A�=�B\��0�5G,��Gc#c����e@�[�c���َm(5$w�����=�e���#X���4��u�2AmH��"#z=���J�x;��Ҳ�R@'-;σ���"5
8^���[!�`�(i3R��ak����`T�ҩ�	r^W	��s��G�z��eh��/��A˥�'ܤ",����^�� �YW;C��U���='����{�6�*F=ॵ��@x�� �<F��1�4q������dz����NR�p�+yG_��\�R�n�G-������+X��FJ���-x�l���ɭ�&gQ�</Sn��/Tu����(�	���s�}�n�H�L)��{TNA���3A�Q���jμ���l�`�g �@�VҒm�HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍz#' ����u��f���`_���pR�_���0����Max��9m3�4��L�O]'\gWg��	�Z�kfc?�#	*]]�iI9�o«IX0F�M��&Y��V�����^����Iy���n���"sS<�0�zG�������&G��+�t2�����V���V�%�1�E���!�nb_X�XV�b�z'hۉ)��d�7�qĘV�52SG�U��@at3Y��P4��7���E�g�������(ӈ���m�r����7�wtMM���j�=Nb����d��i�8���nF���<�W�.�P�	��
�Q�}~�vE�s}�US?�a\�L�O�c���l��,+dN�<@Iv��nt=:��:5A��p/w1z��ӊx�D�Re|����x�.�<������{_8�Y��=�}�Vݨ��}Dq�f�S竚��ٓ�D�=����!o�_"���1�K7͍��|��W&":�ݚ�Н��V��G !]�~F��Ai)̿��n������//�ƍ2���l�~�vE�s?�s^��ɷ��e�ݭ�]�Z�o�)P<�ܓ�Y�q�9�ͭhy�`�w��v1a{J��*:k(v�x����E2b�z'hۉ)��d�7�q�L��@�a��FD>�v��Pn<���@���(9[E�g�������(ӈ���m�r����w Xy�FZ?=��X��/�� �m�Ej�@���(9[��nF���<�W�.�P�	��
�Q�}��k�C�-�+�g�>U�CC����눸�)IdN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H�����Yu���*Y��b"Wfי�b����{�6�o� c ���)΃��_�mS8<�n�ݚ�Н�t�R!ME��ߦ?�~F��C~/*�$�*�]�`u����p�5�"��[�B���p�8����Q����.��$���g�e�㫷%�N���v�9�ʘV�52SG�U��@at3Y��P4��7����*�R���Amr��8On9�*�����C.�u�X��I�ՠ�w�O����;��O�"��H���~�����l���X�� QT��0+��?�A���9-��4�1tSjv�!�`�(i3af��pD�Ї�6~��ȓ�FG����^E4+у��b�Bϱ�����ס�07Syv�Jы�^�)�:5A��p�Ra])n#���r������.J7h����ly�P�r��n�Ŀh$�*�]�`u����p��8��V\�J#�	g��!�w(�y?
�:qEp�;�P�t�5!�`�(i3�V��G !]�~F��Ai)̿��n��_�R��U��@atA�ᴽ�xK���&T!�`�(i3v���,Ͽ�2[QvA�%ρ��r�}6�/S� 8��/��u@hy�`�w��v1a{J�xF0�Ņ��k��M���k�C�-�<�ao���CC����.�<�����v���,Ͽ�2[QvA�t�G�+,�!�`�(i3�5ߧE4��!�`�(i3e<�Ia��lb~*��s�&aD�4�X�X�[RP� .���-a�˩��'����u��r���#�-�p�~�Y���Wql���8z8�t�RL�	��*����Y�U���f�6l�}sf�e�}s�dKa���^�uPϿ.U�d�#�b8�Z���f!�`�(i3�V��G F��x�⢄1@aw5�o;z�j�ĭ�=2�������4�T��Qm�5���J>ni������Cj����tL
�8�[b\!�`�(i3CQ3�u�(���!G�{s��?������xNet&�U��f�!�`�(i3uD�*';;���41IL����֟D@��[����F}���V6�9�leD���>E�%��*d��:=�;]C��ZH&R!�`�(i31���~!�`�(i3af��pD�Ї�6~��Ȕж�{�7�	��*����Y�U��3Y��P4�|�OAn�!�`�(i3��Ě�����}Dq�f�~�vE�s?�s^��ɷ��e��������A�V��G !]�~F��A8z8�t�RL��}Dq�f���k�C�-�+�g�>U6���z�S�D����P"G�wk��%�])�+�[��m�U#��Э�@�:5A��pw Xy�FZ?���3���α� �m�Ej��m#?����W�W[��m�U���_R�ݚ�Н����F��O�!�`�(i3�;b�-�2��;�P�t�5W?�;�끣�os�鮊��~TX��7Ɨm�zD���'$3���WS��0+��?�A���99<���F�8���U��@at3Y��P4O�˰�]qv���,Ͽ�2[QvA���x��~��Y &���B��2�k1�h�H��*��s��R�-��J!Ҍ5`��/��kOT�V��G !]�~F��A8z8�t�RL�h��N�M��z3:��K�z{�� ��C~/*��f� .):�@��A���k]m���݀γ��du����p�����+X��FJ���-Yk��P(I��MV�,oy4k���Z!ƍ2���l�R��ak����`T1�h�H��*%�줝v)ڥ����Ⱦzk����G7```+�8z8�t�RL��%�.�E
�ߦ?�~F��C~/*���2�*#M����ge�`���*1��&g�hh\�F�u��� �<�5Ɂ7����W�W}c��ko#ƌ0Q_,�8���U��@atA�ᴽ����rv:�F!��D�����q���<�W�.�P�	��
�Q�}t�,�NL}�="��x8I�t�2�q㬑^)�G�B�+�WdM4@����[y�K��z3:��(���!G�{s��?�����T���E����X��O���r����!�`�(i3!�`�(i3�>=���#F}���V6���w�?�R��y	����F��،�W[����Z�,��#�2
��e�������m[�LEE�S�A@����d��-��!���Bvy˥�'ܤ",��Gc#�����O�m���Ar)���r����!�`�(i3!�`�(i33��0��e��0�U+�qbp@��x�bG�Uew���m�|����x���f�����&Sq�a;Uйc�e�ʥҔFܽ���ly�P�r��n�ĿhxK���&T���sK4�֢��s�KȔж�{�7o9c��@��@R�^���!o=��MYwO];;���41IL����֟D���Ef���@8:�"�Nec���P�ߚ�6���'HY-��
�C��n�%GPM�^-q�x�l��1:�N�*�x¥������]n��-��%{.�V#?p�&���A	{K�tU�P!�`�(i3�gCu(o?C!�`�(i3zR��_��m��3��p���H����Q#�?���;���Nxk�~̔=Z!�`�(i3^P��:w0I� X�1�;LV^Š�r��Lo�_!�`�(i3�2*Q=F�k�mD#V��A��`-2Y��kک�x����y���ݫ�ф���F�)�_�������� "5�]�B�'��a�F�,�U6�Q�L���/��@��:$����z�����	�;�ݚ�Н���"����M몴PBoT�ݚ�Н���_(x��`g�%Y��̗0z�cUL��s@OĪkew���m�|����x�hH�
$;�?V��j�c�;J�*%n�d��}U؄�k]m�����2�¤Z���wj��89����X�G[��O�Z�_�m��+�Z����y�MC���d��R�7h�,b0V�u�Q�ݚ�Н��
�I�>y!�`�(i3�U���A��y	����F��،�k�+9=���-/E8�)�[���6�X;p`��L�溥����v�8:��|`��'J�	�LÆ�c�9ʼ��$$o#[�L\��@1z�+J���5���Adu�5k
��Fɴ|�O�j�gh�䊉��	��J�6p�N��2��,Wc��I$��:�e�h�Ϧ^c!�6 �ef�&�2�������ȍry��	Y��
�iCTl�������l6���0�&�ͭ�U젩`#�4>?� �1��ɕ�eY�����w6YmC,igu?V��j�c�
���!8Z鎬�������(����,F(dA�F�u����ӕ�![���ݚ�Н�p�n�����^����+�g�>U�#!���e����M���^����Hb�2�Ǐ�t*�����b�氦�=��X��/{A�dha#4�8�e
��'�i�*ڶ�UKs,��l�?�C�gXk>!t�7ń��,�HK�n�Jt�gc��u���rQ��qD���Hb�2�Ǐ�iA'R�	��)���sf�e�}s�dKa���^�uPϿ.U�d�#�b��R=y�t+�_0c ۘ�C�r�s=��X��/�}VV��5l+��@-�-'͏������ӳ3z�]��t�iZ]XF�hx��G��!�`�(i3U��֜��3!�`�(i3X�PC!v�@[�JJ1��P�M��,���9^-���.��֞�������i�4��%�;��g��cH�wA�?�W��7E��n���8��T�h���}둮j\����C$L$E�͆عE���ؼ(�K�^��Q��G�S>\.�!::tm�0�i.�9gh�䊉�䞘gx�n�W�����v����?�dv��oTN֢&@��&�_F�k-��苇��Fe#OOJd֯��|��p��PIQ#�C,0�?��ʉ��%>�rG��M����{����"�2��}��CϾH�)v���,Ͽ�2[QvA����D/@�2��}���zgm##�v���,Ͽ�2[QvA�gN|���!|Z���wj��89����Y#ѥhB�@o��[^�}� u��=��5W_����L�,\ަ�It��+g[�N����p$��<
DN͗&8�,�8��!��L�E��w*��ܙw�F�ݚ�Н�rM�e<�!�`�(i36�X��U�o̥�0�L�p~z�r,,���9^-�ΡKCh��(	�G��^����K�7����&Y��V�ǣ©��$��:�e�hfH'��!�i����VZDf�?ǉ�=�O�G?X2�K��2WI'�=��yp����nZ���t��˳3[�u8��M�g����H��bf�?ǉ�=̇i�d�?�4�0 L?�p���@Z�6[��u�9k�\,���m�
��,!q�\E��0Z��0�Yǆn�Jt�gc��u����ժ*)xJeq�\E��0�>���W�n�Jt�g�v1a{J��OSu����І�TI6j�"Hs`]��ä�l!�$�"��`� �3�<����,�ǰ&k��������a5���֓��@ee��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcM"o�N. X��(��n��	�(��N�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�B1����!�`�(i3�U�s
ƺw4�f/���l�l"��l䋬5Kq�1@��b�tS�SaqZXr&ߜ�>�]�P8�.�I�A��ht��p�éR��5�"��+�������B['u�_�#g� |���R(!|���fw;k<A����'�QDn4��F�(=2�F?�\��Ih�	�;B�"�ɚ&����'�h�5,Wlr�r%)cAQ17�b�����d���!i���jSA n2ϒ���=��pȠ��ղ]��G��-y�� ����i9vo��ob$fAԢ�a\�\���V#��p~z�r,)����2 ����i9v��խd�g��;�!�`�(i3!�`�(i3!�`�(i3]q>�A�	?�t�ϗ;��|B~����`cg��L�*� )�\�~xy��Q�^e�H�qfP�����5�����0��+�!@�N����f0� ���S��B�xL�����ܢ��i������^�
8�.�O��QK;ybl��Tx�^ʩ�}���2�4帎}~�K��8l�=9��ŏC���-�o{s���CQ�����m��I!EE�f�g`�KU��9��̵����V�@1M�"��b���R��r܁8�7�62'~3\�]�0�
n�f���=��YV�g��L�*� )�\�~xy��~�_1�H�M�;����'�̗�����AJy/���K�4��L�FZ�1����ǲ]��Y�@L���d���!i���jSA n2ϒ���=��pȠ��ղ]��G��-y�� ����i9vo��ob$fAԢ�a\�\���V#��p~z�r,+������Π��yGb�s�-xe1{�;���N1v�0=i�R�c4!`�d>�c�n��N.�6�����k$ !�`�(i3!�`�(i39�O��F���{S'������,�ǰ���!�Ab�f�s�GB�"�ɚ&��f-m�b�,�W7�_��kv޶GlR�c4!`��0]A��~˼��H����8����F)�~��[t�Y813bQ=�3�� �֤D�A����<g�?�d���&�_��5��0$$��
�5L��m}I>3d?��������G�9I��@��~��q6g�yF}���V6���0�] �v"��%��+V�R�c4!`�d>�c�n��N.�6�����k$ !�`�(i3!�`�(i39�O��F���{S'������,�ǰ���!�Ab�f�s�GB�"�ɚ&��
$hu�x��j+����@~H��k]m��E�M�����x����~mW3E�-).^QQ<7����ͼAԢ�a\���y>'MM귈nIg�RJxo>��-�ļަ��P�5��/dV��H(�T�O��{Tɀ�$����nQ�rVA�H��%�'{}yw~�귈nIg�R,n��N�d&�.�_�L[� �h���Y�CR����]#��t�ѕ1��ŦLZ��Ѡ��>0�1ۍ�h �=�)��=���!�`�(i3!�`�(i3!�`�(i3}Y;�jn��9��稕/Tu�����_&���*���)ei��h��N�M��G��-y�� ����i9v�A=K�����_
�u�}���:D�_�k�Æ��%N��� �"�W�A�&hH\�LZ:�\�Ԋ�{Tɀ�$����nQ�rV~��s�N�h�5,Wlr�r%)cA�F��=��g�]@n_���?3ֳ���[HDȚ��wz;�|�����I�HM���#g��I�mV�Z9I��@������Z>��~��l������IV���@�\#��hvl��9�h �=���_��')�c�n�RÆ��%N��ݚ�Н�!�`�(i3!�`�(i3!�`�(i3}Y;�jn��9��稕/Tu�����_&����=/����6�h��N�M��G��-y�� ����i9v�A=K�����_
�u�}���:D�_�k�Æ��%N��� �"�W�A�&hH\)�s!��3�귈nIg�R�5��/dV�L�溥����v�8:ۛ@W:���#���F��*{�욋�Օ��qvdЧ^{�jЅ�l�H�g��cH�wA�?�aHǮ����_G3w�
|:
@�!]�݃��x��q-��#N��]#��t�ѕ1��ŦL�_���`����Fp7�D�_�k�W�A�&hH\�#n��f�-�o%�_�*�@W!�`�(i3!�`�(i3!�`�(i3!�`�(i3V[B�5�m�x���|��\� C&����q��Z��2Q�g)/<�C,�#�ݗƩ�@�Af8�ٕ��(�W�!Ċ&���X�G[��4
� �b%m�Y$� 1 �ټ���\� C&����q��Z���J��"���p
v�ݗƩ�@�Af8�ٕ��(�W�!Ċ&���X�G[�D��$	�%m�Y$� 1\�]z�+����3���΢#�7�
���?���A릂4����af�G���Fri�u�q��k�ʆ-�̍;��!?j?�d���&�f ��˥�'ܤ",����^�� �YW;C�ͼ��O���M�{�|L���u��y�ڭB��2�k1�h�H��*F7	G�<�*��s��ꮂ�n��;��f���-A�¤�x.�Knq���;W��ZLN�	����n݁Fri�u�q��k�ʆ-�pd�
���M��7��(�JZ�Vk�;��|B[���ɐ��5?�&P-ߕ�L:�,�����^�� �#���f��n�Jt�g���E�*��p�O2!?����^�� !
=�vv�>&KӔ�o�J���" (�P@L0��U,�W�8"M�5�O�%E#PR��ak����`T�ҩ�	r)��f�� ����7�|ʔ۫;��w�R���y�T$����FD>�v�ހ�mcQ���+O*F=ॵ���:���K���~N|e���b�!�`�(i3�h��N�M��~��f�!���zՠ�~��q6g�yF}���V6M��C��]��ġ��,�����Q®��zՠ�����Z>��~��l����r����!�`�(i3}Y;�jnc�n��`�7�,��n6�o8:4�I���c�90��G��6�iI9�o«IX0F�M�H{���<�e��BFbs��2[�a��o���H�RtV�^+���G����$�\%e��}Dq�f�#� �,W���Ǉ�y!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^e<�Ia��la��o���H�RtV�^i��H�p¢	�B�d���%���Ԝ�}Dq�f�*�9��.���i��/�z��P��*|���%>�rGO�D mWN��Ě���aT��3G�IX0F�M�H{��'�n�2�M�]��P�),�ѕf�f�_T:5�����2������}W`�J$˄���Z��s->m�9V�ZP�����Fz��Ԥ��ht��R����A$�P������5d�������y�:Fa�7�����~�Lk݁ 1���tw�i�Չ@�^��1���"sS<�0�zG�������&G�/��@��t��ܜ�[�dN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H�����Yu�������&G!�`�(i3͜��!?@K}�1U��VP�CXm������>?��"X��[��0�����J��sr�l���ԵU{fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx���Db^<�..�4��<qs��aT��3G?�d���&��ٸs3}A��O�����N���Pm���֛�l����c�n�RW�A�&hH\+��O�r!�J��:����͜��!?@KE�g�������C�tpYx�J��sr�l``�^��c����,�ǰTm�v��G�3��P$���V�6�/�@޼�	�f�]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7�p���"Z�v��!\���F�`yx�>�+X�M?��y��#�-�p�
�p�	%6!�`�(i3!�`�(i3!�`�(i3�q9+t�}�;b�-�2�Nh���W<˥�'ܤ",^� ��B!�`�(i3x����E2b�z'hۉ)��d�7�q��6[��u����@~H��k]m��Z��h%�o7!�`�(i3E�g�������(ӈ���m�r����%��C���Q׆��p0�Ĝ(�IyI4.Y�fV�l!�`�(i3��nF���<�W�.�P�	��
�Q�}�L�����B��2�k1�h�H��*F7	G�<�*�P�ߚ�6�h��,���fR�,� �GR��shbvk~�#x ��M��.ᬵy����uq!\H�q���3��`��R�`�mQ�x�z�oi���:�R��_k�s��c�7�wtMM�0�5G,��Gc#�����0o� c �,��m�ܻ��_
�u���nk+ߜ�*�l8�b(������l__�I����J��.��c��D��_�W�.��;�#��&�qҸ�2Mz`���^��D�Ϝ�}Dq�f�q���3��`��R�`��ƍ ��_~�:N�����;q�{_8�Y��=�}�Vݨ��}Dq�f�q���3��`��R�`K��"��zigzA=v)����;q�{_8�Y��=�}�Vݨ��}Dq�f�R��ak����`T�ҩ�	r�MBD��������;q�{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^e<�Ia��la��o���H�RtV�^��~Щ�!�`�(i3!�`�(i3��X�z`ʙ�SQ��?D�8���6[��u����@~H��k]m��l��'�cv�A�
^^3�V�C��k���a�K�v�A�
^^3�V�C��k���T�7:ܑ��y���8���/��R�E����Q׆��p0�Ĝ(�IyIC7+h�6u�!�`�(i3v�A�
^^3�V�C��k�HvL)��9�;�0�*:Wfי�b��}!D̅����<!GO#(��cS�c�X�X�>c�.A�x���0��"X��[b�&�,���Nh���W<˥�'ܤ",�����D�-)�_�S��R
�:qEpNh���W<˥�'ܤ",Ц�} m���o8��l�x����b�'Be��/=��v�A�
^^3�V�C��k�HvL)��(o�ܷ��a(􆿳�pr͚]j�Wfי�b��}!D̅�������.�']u4c!��mJ�0�6���+�t2�����dz����NR�p������jp��X�z@�Af8�ٕ��(�Wa�su�I�q���3��`��R�`��ƍ ��_w�?��g��U-�ew{�I���0�5G,��Gc#�����0荛y�(*N
����\� C&����q��Z�����gf�r��}�%DܭD��_�W�.��;�#�A�=�B\��0�5G,��Gc#c����e@�b�������Cҷ��ep"�ߏ׍�B��2�k1�h�H��*��\R�ݚ�Н�Z�,��#�2
��e�������m[�X���2:#eh��/��A˥�'ܤ",����^�� �YW;C��U���='����{�6�*F=ॵ��@xݵ�Q�n��T�\ ��;��'yJ�V�C��k����?dq���z����7t6>�&Չ��%>�rGO�D mWN�s�Yls��8��GM��i��.l�x����b�'Be��!PɏPv�A�
^^3�V�C��k�HvL)��6�5Y�S;����1H}�ɐ��/�Æ��%N����[����2+m��h�����H���ʖ��	�_C*ζ�I����;��P�jcd�LO����K���Yb�Y>�fW�N
%�Rk��4��J^�B^�����f�L��'��UCmV��!jG};�;X�ӛUi]�g�^����H����q���3��`��R�`�mQ�x�z�oi���:�� �y鎣�N���!�`�(i3u����p�����+X��FJ���-],��%s���@����^��C�=�g4�B��2�k1�h�H��*F7	G�<�*J�QF�n)�>������$f��_Ub�F�S�1 ����F��O��|#HK��=�O�-v�*�Va�irv�A�
^^3�V�C��k�HvL)��E��PT�Q׆��p0�Ĝ(�IyI�1������FZ�����J�d�@q�2������}�G����_�mS8<�n�*�p9��n8q����ij\xD�Z�=`|;&o�f��ʭ.��;�#k�����a-����|K�-oF{��=��,��0�Q�-�3P��H����^���	��L�� �[cz1�� ���@A>�0T|��h�؀!�`�(i3�e��	�K�D��_�W�.��;�#��&�qҸ�2Mz`��Q�kŕ��QH�RtV�^N
����\� C&����q��Z���2%�ɛ'�F7�GhsGS��c��0�5G,��Gc#�����0o� c �Lʳ�nsR����%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��j0C.�>��V3o�Ik$	S�uimK�ֶ����6�o8:4�I���c�90��G��6�iI9�o«IX0F�MR�c4!`{ਃ�6�����"sS<�0�zG�������&G·���~X� ����i9v^�?�K7͍��|��W&":hDJ��3�D厺��+�̟�1dN�<@Iv��nt=:�$r�t�}ik+Q�h'�Ȝx�5W ��̫(� h�ҩ�y�}�6f&rG��Hb� h�ҩ�-|��Y�$,K�9+�/���p���Ӗ���������5����u�h1�M?��y�!�`�(i3�m�n���Y�j�`M�4d	t�`�I��W�T�TN�����%>�rGO�D mWN;�jmT�#Qw�$��Z��/�dW���3����V$=�b�oj�+p�K�J�iN�S�"�����<om����=&%'�Du��r��d�tu����a{���Bf���oj�+p�K�J�iN�S�ԝy'��Ra])n#���r����>�Q�c6�����-ќvlr�{��|e��0�U+�qbp@�!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�MR�c4!`��]��R�3S;nc,Ec'�\Y-φ��<�6�@a� ��fFMqlg{y����i�q,?5q��7���9��e���W� �{Z+��r$ɓǃl[�Ƶ�1tSjv����q�D�i1.��2�8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩ�y�}�6f&rG��Hb� h�ҩ����q�D�(�Ha׮�#K���~N|O`�� \)���F��O�}�	76�&�� Ӗ�t$�)�vx��SJ��2���P��*|�t����k8�J��sr�l���t�T��?E-h��`f���sd�G}%����3f闶P���`�3ޕ �7�癆cgQw�c4~Nr_�mS8<�nt�{#	�x��J��sr�lE�g�������(ӈ���m�r����*qA����6\�4�@�� �-j�1tSjv��
�t��T&���LQ�/81tSjv��H�����S>4�mDWQ�g��	�0�=<MW�-}�	mp :H��\�P/0G�D����M��p�#���F�Q���*���-����!�`�(i3�4�	���+4��8��q����A��>��������w�w:�!�`�(i3�j���%��Z�H��q�e��0�U+�qbp@�!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�Mcny��&�M��xx x �i�{���w��k�����T�}ɻY~�y�����[�T���Ӫ!�J��:�����#}�{��9�2�LK7͍��|��W&":��;_��8W�w��fD�]C�1�vv8��
�1�c�{����@&^�T ����Օ��qvdЧ^{�jM|�"D5�O�%E#P��C\��~g��tcb�A���t�T��?E-h��`f���s����a���s�*�I��&����!���� Ev�P"G�wk�١��	;q}u6��\����m��3��p���H���F`���G���Cҷ��e�ˇ�h��<�W�.�P�	��
�Q�}N}�m��{t<�J`�) �U.�\�/bғ�vq�\[$Q��
�̞��>�h�5,Wlr�r%)cA�z���a�1;Z�减u��>���e��0�U+�qbp@�����a���'���_�)���p��b��x��f��]�!��	Ǹ�y85������GyV���2a� �������!�`�(i3�ˇ�h��<�W�.�P�	��
�Q�}{y����i�q,?5q��7���9��e���W� �{Z+����"sS<�0�zG�������&G��+�t2��&����!���� Ev�dN�<@Iv��nt=:��:5A��p�/��mS%�U.�\�/b�}�Ш���my$�N��o�/���;�B�'��a���p��b��x��f�dN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H�����Yu�������&G!�`�(i3�#}�{��~v� 1����_k��iK�0z�cUL8�l�#���P\�C�Lz#��#�'��o�u:��_xۏ�:��"�#}�{��~v� 1����}Dq�f�pT/�GS�)���܇�b~*��s�͝������̟�1��H(�T�O��{Tɀ�"'��&އ��-/a8!�`�(i3M*KJJ�[�4br����&r��*u!/��"���,Vr!�`�(i3��:e ���N�R���Va�ir���e�T���U�._��L�溥����v�8:?�'����-����!�`�(i3�)�z4J����aGl��ˇ�h��<�W�.�P�	��
�Q�}!�`�(i3]���-_!Q�U.�\�/bǴc�1�RG�p�P�m������� h�ҩ�!�`�(i3�YN
��)ehc�f����YN
��)en�@��BT��}Dq�f�՝� s�#���k$ !�`�(i3�YN
��)ehc�f����{_8�Y��=�}�Vݨ��}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j �_�ȇLШ��+����-Q�OP����,�ǰ����adp��e���W���e����VU�簦��E.t�