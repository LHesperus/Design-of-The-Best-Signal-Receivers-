`timescale 1ns / 1ps
/////////////////////////////////////////////////////////////////////////////////
// �ļ����ԣ�		ģ���ļ�
// �ļ����ܣ�		ʱ���źŲ���
// ��˾: 			�Ϻ���־ͨ�ż������޹�˾
// ����ʦ: 	   		XLX
// ��������:        2010��12��25�� 
// ģ����:    		TIME_BASE 
// ��Ŀ��:   		MultiFunctionSignalSource
// Ŀ������: 		EP2S60F484C4ES
// ���߰汾:  		QII7.0
// ����汾��		V1.1
// �����ע: 
/////////////////////////////////////////////////////////////////////////////////

module TIME_BASE
(    
	clock,
	reset,				
	PROG_INT, 			
	INT_ENABLE              		
);
//////////////////////////////////////////////////////////////////////////////////
//�������IO���Ŷ���//
//////////////////////////////////////////////////////////////////////////////////
input									clock;
input									reset;
input	[31:0]							PROG_INT;					//�����жϲ�ѯ����
output	reg								INT_ENABLE;					//�ж�ʹ���ź����

//////////////////////////////////////////////////////////////////////////////////
//�źű�������//
//////////////////////////////////////////////////////////////////////////////////
reg		[31:0]							CNT_FOR_INT;

/*********************************************************************************/
/************************************����ο�ʼ***********************************/
/*********************************************************************************/

///////////////////////////////////////////////////////////////////////////////////
//����INT_ENABLE�ź�//
///////////////////////////////////////////////////////////////////////////////////
	always @(posedge clock)
begin
	if(reset==1'b1)
		begin
			CNT_FOR_INT 	<= 0;
			INT_ENABLE		<= 1'b0;
		end
	else
		begin
			if(CNT_FOR_INT==0)
				begin
					CNT_FOR_INT 	<= PROG_INT;
					INT_ENABLE		<= 1'b1;
				end
			else
				begin
					CNT_FOR_INT 	<= CNT_FOR_INT - 1;
					INT_ENABLE		<= 1'b0;
				end
		end
end		
/*********************************************************************************/
/************************************����ν���***********************************/
/*********************************************************************************/
endmodule