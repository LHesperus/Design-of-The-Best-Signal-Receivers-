��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G0��@h ���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����pn�R��}"C��dKBE7\F���r����&$9g8�M>PFWD#�z":���ӳ��_�x�$t�`a\�R�F*}Ø���K�ZF��W��`k�ZV"���:��#tC������s��n�
8JA͎��T�k� ��d�n}K-J��K��z������3�z�ω���D���+��ԟ���F72��{L�8br�.�/�d�������4�;���u�$|�>I��4�Y�YrT�#ϯ��=K�)yH�I@'�ew2�\�蝆�u����l�|���j>�9�	)�ň��h���N�$����/pZ
OC`��<�H6i,ER��DT*����@X�j,Zs��?��n;�|-���g]��~����B����Ls�Fޣ�@�ѥ���vH,�uS��wQx�vyPTa�������N�s��< 
��݇� U���/8f���p�ny�(�[x;-����o�I\\+�K�&�a��|����W�%�э�j��~o��;��|Bm����ܸNɇ��nC1�,n���&���N������8��U�
ث*����Vs���,��}�_��x�j؀O��u�>�����j�3��w���j������x��(���a���<5(N����7W-��L�@�y����L
�T�p r��|���-&�TfH8E^���G�38���E�x��_���|5�$Ծ蒚�(
�ݐ�s)9l��(��^�mD>�0aH%f���eϥ�2@��9���Ih����M�nGpԆ\A&���F�\�e�}˪�ckx��6֏�c �l��0u���ߏ�e�e�PkѶ���� ��.*�_n�2�HG@����)��>]�Լ�c��l��e�E�s;��Ӓ�T���W�W��Y���^2�i��E�V���Z'�YQd#�;�Z��`�+N*t�����,-�qĬ�z??��'�`7���X�ͮSN,Sh���$�(�+��M�.�.ni��l|al�g�Bp!!v*!��x+���1��Lj�XW=�`H8���;��pmf����K���$��%�`�ny�;�ns)��E�$+�>����]�4��z�tx������89f�ԝ�f�Q$�9og�`�b���z����j�V��v�g���rz�\�2��s�#�<����X��|�E��Ց�x]t����Z��+�>����)�i�~4���Z��_"����$�Zj�V��v�Sw��ꆚ�>����9�H�o����8�!�r���=�T�����0��GB7 Q�s֞f�4��r���7��ӫ�Wt����֤R�g�(0e���؝�Nu��궂Oho��]F����M�m>OM�Ѫo���>�'�f!���ٗ�U-f B���R��#�Ulg�69��1��`�+N#�H��h�3#ب�Re���L���$��fF�:ަ�:!�?�)�H�vƖ�"k@:G��ؠ��E��9��-K���}0x;E8�I@3U��9��q�b蔹Ci+�/0�?D5=��<}ϼ 8�����1mS�Q�ME�EgJA��3� ��w?����9�b��A�����w�6����5B`���YK͊+�[�q���ff�u��T;��n��&�;����H�3�s�3*]�yRy��BY�/�����	�d*k�u`�E��a�"�u;�:B�@�zO�üx��!.�R�9�I�1�\�^6�샺���j���Jm�W�(�P�Ϣ�X�b�T(yL��탧m�$�8��!��8���G����7�Q���==�^���@Z��hf�.�?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��r�����A�F�7���3�GXS����E@��~���($�J.���
2,w���~�?|�[_wȵ�e�kY��Y+]��=W�֯��i@F�5�=h�GD�#�̔"v��ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l�������+rb��@���,������0��D��L���_�L�3��0I}.��dPc)y��0��r2�􉢔�S�����5W/�؏�<
DN��E����F�Z�>)��p40�zɈ4X"��D�����ˇ%Ah�%4
>��XP��������kV�^�o�\9a|�����#�ڊ<?@Pʶ=������Y�}�f�����g��������\�vňu�,�s�K��U�DG�p�P�`�>:8�A�/���a
%���A�+0�l�R<�Q�(*w��k/�z�xEQ!�`�(i3v�ј�"��Z鎬�����X���*�V��*J !�`�(i3��|g�Y�'���Xw�,bxqX�2�����Vc�@�Q�3������o���g��m�wR)$�Cb���ٜ�]!�`�(i3v�ј�"��Z鎬�������(���	t�����"j���b7|#9���EOJ�uxm�5���u�L�Y%T��BPe.��xu	���S8�P䴰^MW� ���t��!Z`x-���ˇ����#oMZ�n��[��{_8�Y��=�}�Vݨ��E�d��",oMG~�Յ$�O&�c��Et��q���U�+Ќn'I�+��x�v/csO�LYw9����-��%Mό���.Ӂ��̰�!�Xy|�W�E����F7G#+��\w��0]C�4M/�S��ݡ��1��Y%T��BPe.��xu	���S8�bM� 2)G��8���/��,bxqX�2�����Vc�@�Q�3�y=/i�Js���7`�gnk� Ɓ����[;�W�@���+g^l����^����>4�q��]���>����C�x�j؀O��w���B}Yl���#�]�!����M[��Ǣ�\�2��s��+�w>���]2�y�Z鎬�������(���	t�����"j���b7|#9���T#�3�["����:� %Z�P�c@IE�U����S8�P䴰^MW� ���t��!Z`x-���ˇ����#oM|#9���T#�3�["�Yr/r����
y��@IE�U����S8�bM� 2)G��8���/��.aX�bAKj�V��v`S��|��ɕ�(�
t�ژq���U���V9{)=�?��3�;T?΁)��TD��(0̈��N�2e�5�ONG2�꺆���$�@O�x�7�k�ZV"���:��#tC������s��n�
8JA��C�Y�)��NË�����8��z{��E�EYZ/�矘��-n��I�?g�f���\X�<����8��UWJ��)�-�nC/$�m��P��I��'������[��CCLn��S�W#w���	(���B�� ��I�=M�^"4/���^���4"�ND�A���@�k��V�4���|;��7����'���ɋ��9�?m��W�m�ꭂ?M6����)��d�j�	�b!��u��K�&�a�nS�dB�^�vtiDL��Oއ�?t},�׉é(.V�����ҟw���Z9�+	�xg`�H�4��`t�A~�@����gG��s 1!m�vIN�E����FZ鎬������_�,��T:���V�T���!�`�(i3�d�٣���N N�S���DP֞ ���U�B�r���n`5�fK�\w��0]b!��uፆJ�g�*�~������+�J���q���U��@����gGm��s&}o�~��w3*)�g��OZ鎬�������(���/��A����d�a�4$�b!��uፄ\�2��s������x~>���������q���U��@����gGm��s&}o��b��M��`M��
Z鎬������_�,�� ʔ.te`�\1^O� �Xz����d�٣���N N�S���g#j�V��vt}���#��n`5�fK�\w��0]b!��uፄ\�2��s���1�, �_�S�
ut�q���U��@����gGm��s&}o>&S�XQ�?㐌�PB�Z鎬������_�,�[/�cWM���Xy|�W��Υ�d[g�d�٣���N N�S���c��:KYЙMǿI?��t?�@��n`5�fK�\w��0]b!��u��K�&�a������ +���+�J���q���U��@����gG9��I+nXB���2#�E����FZ鎬�����
!-�n[�=�5x��$*���!�`�(i3зq8�Ј'���Xw�j�7���5�%]���a(􆿳���2����.��DP֞ ��+�?�!�`�(i3�E����FZ鎬�������(���Jם����"X��[��Q[R�7����n9���8��Ս!P����"�,�>E���]�!����w�Հ�[�=�5x��,����I�''Tq�q�зq8�Ј'���Xw���,D�>: �.��B<�L�V_!�`�(i3��Q]� _ό���.�}�
�?����'�u�Wql���8�{�����7s�9���o��S8��y�)xʔ���6��	���`y����@����gG�F��o�F�M��:�j!�`�(i3�n`5�fK�\w��0]b!��uፇ,��7-u��Y�r!�`�(i3�d�٣���N N�S��+\�g����)e�������:y����Z鎬������_�,�n�j�<�� �e�d���e�Tnee]���+�J���q���U��@����gG�F��o�F�M��:�juҩ�6�f;�n`5�fK�\w��0]b!��u��c�r%��'L"*!�`�(i3�d�٣��c�A�L'���W	ܷ�4D�P��dq�8���/����,DU�m#j[��NۥUn�.�k� ����Q]� _�rs�i�76b�*ҒT"h�p����t%��zxa(􆿳���2����.��DP֞ �'��L�������:y����Z鎬�������(���:���U��^"4/���°������R�wX��}�
�?���v�)y�Eh�ѮYț!�`�(i3±�sR�{F�(R�?j�����B{�J�q޼UR��-r��|ڑ�8�
,FI�}�
�?���^(C<�@Km��}!�`�(i3±�sR�{F�(R�?b02�O+c�FP_4D��ɍ��зq8�Ј'���Xw�j�7��a(􆿳���2����.b��1pO�/B��͵h.?�al��E����FZ鎬����;��0��t4�6@|����h[,ώ ���]qLM�!��T	ܷ�4D�P�>�s�,�H;��|B#��7N��%�эȈ]Z��������;q��b+}y[��+g^l��+��\���E�`JcU�q9+t�}�����~�A�qIp��K�ڶ|e��DE(_
/�Ƀ�?PA�b�'�wJ:^	QW�Q!r�{F��#�����R.P}>C��<�j��۳a'[��%�э�X6و�cµ�Je��v�i�:`�+P
��K���7�`K~��'l/7w|]P���V�-��&�t.�}7�`K~���?g�j�P�񭩶��&�t.�}[��N���ҟw����f�\%�,�F��P^��"�م2�w����r%�4¼�kF*�L��!�`�(i3!�`�(i3!�`�(i3���.ݍ|��C�t�ؒ�9��t`�<�C,�#aT��3G?�d���&��v�<���+�+\���;TŬ���IY����[e0�~�zR4 :��	��԰/�&7?�d���&�N-Y&yo�qS竚��ٓ�+�Lr·���Dhƀ�^
�����|��*ȑs;��|B���r��������n9�u�#�$IX9yAjq2w���P��vZU2h�d�+�q�Q`����"X��[��Q[R�7d=��¾ȼ��.J7h��F�z�>�/~�[��ϸ�"^�j�h�5��
�YW�S7�.�,\����g�T��ο�^"4/���6�-��ӸT"h�p����8.����6��F��8!�`�(i3!�`�(i3!�`�(i3!�`�(i3im�x�����Z���ot5^ݿ牴)e���Ô+;��2ќs\5 ����.��?��wO��Н�:���M��:�j��G慧1���~!�`�(i3!�`�(i3پ[���-[�g�DPp�Q� �_tta��������G��L�1p/-��9mh��n��V�%�16�����uD�*'�xѴ��>3d?���2��HO���u�#�$IX��ݣ_-�iJ5a��!�`�(i3!�`�(i3!�`�(i3�_��U&���8��Ս9�y�ł?V�fc$��b��X���&R�n��Zn���EU.�(���[0RCm���Ӱ�e�����U|�W��eg?��v9���r����!�`�(i3!�`�(i3Q� ~��HN��R��?�d���&�af��pD��8�WI�AdS竚��ٓWqo
jk��P:�z��������*s��$�Z;��|B���r��������n9�u�#�$IX9yAjq2w�f���,(���B����V_���07��i:��ê���#oM|#9���O.C���=����t ��A�Y�j<�i|nơlП���}��%v�\��ސ���97��EN҄����T�=�+�#�W��5�t4�͎�R���HC���*,w	����ز��@ȼ��r����!�`�(i3!�`�(i3S`�@���=����t0]��2�O2�*�����ϸ�"^�j�h�5��
�YW�S7�.�|ʡi��!�`�(i3!�`�(i39�O��F���{S'��:)!�1%�@YC-�T^*H {��u��]'\gWg��	�Z�kfcM��fZ�d�G}%����3fL����:�YC-�T^*s
9��
���"sS<GYqcHTX�';��#j�ݚ�Н�EOJ�uxm�ސ�����nF���<�W�.�P�	��
�Q�}�߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3oв%u�K�w�c��l�,� ���uZ��_����3Fڸ�>P��=����h���7u׿��� h�ҩ��wӨj]h�u�#�$IX~f�@�f��e��0�UX�Pp42JFf���ސ���6 y2��R�՝� s�#��qX7'��|�;�Ojz�$�AՁ�Va�ir�\�2��s��W��7=#o�]�ʄǑ�+�/Z �ސ���qQ)Ԥ�wԿDomn�MH�Ћ�r�H�RtV�^�2��}���'��L�㜰�� ��'��L��\�b�a!�`�(i3��$���͜ ��A�Y�
���3ʩ�>�X6�j~H�RtV�^�2��}���'��L��˰M{�?I�my$�N��o�/���;!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2�$�)�vx8tܟ}�nEg�N>Z������V��	��y�y�^	#�3 �2r�����~�A�qIp��K������"��2�w�����DO&��Ni�:`�+P�!��+LTQ�g���J���X20�i&<N��M�{�|L�8�YX�s���{
B��T�eq%m ��;՟��}�S�4L_�X:�����f_N��ҟw��
:1�U��������ݚ�Н�!�`�(i3{�d"���ƍ2���lę%��%���y6�T�@�����M6�o8:4ڄ\�2��s����a�v��x�j؀O��@EZ����f�?ǉ�=!�`�(i3!�`�(i3!�`�(i3��.J7h��F�z�>�/��4�y�c�}��w�I2_v��%�<o�;)�yԗKo��1!�`�(i3!�`�(i3!�`�(i3!�`�(i3i�:`�+P��Q���r��Ƀ�?PA,�$$*&�ЙMǿI?UKpm�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�,��7-C_u�y�Ǉ,��7-�P��U�Ƥ�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3��F������0��GP����˚Ň,��7-oc����HL�WUJ�N�������y�:Fa�7������A��Vx���_>
xM�v.���)�D��)�{6�U���.��h_'ЙMǿI?��E��D��ݓ�W���0c���cͧ&U�)j�S�mJ�0�6�!�`�(i3�tU,�Ql�	^���y ��-O$U1tSjv�!�`�(i3�(R\֎u��w�`L�h��=��޵g!�%=F�=!�`�(i3^	QW�Q!r�{F��#��g�+C��s�t}�F��<�����xb�ݚ�Н���F���K�&�a�M����*��q9+t�}�ݚ�Н���F��=�?��3�M����*�'�^�����ݚ�Н���w�w:�!�`�(i3^	QW�Q!r�\1^O� �Xz���%��v��!�`�(i3^	QW�Q!r�{F��#��g�+C��sJ�A7���ݚ�Н��H�����,��7-oc����H�}��ɣ#o�]�ʄ����n�0R�0�iN�
_��f�8
��$����թT��6�F���N�DNl��O	S��Gu��r��!�`�(i3�%t̓�@���{
Bk	䶙%��򴶽!!�`�(i3��+g^l���b��M�-��h���?D�8��!�`�(i31���~!�`�(i3(@X~�H:��}�S�74/������.ݍ|�!�`�(i3��F���K�&�a��i
�i�w)P<�ܓ�Y!�`�(i3$f��_Ub�F�S�1 �fĉ>99��A0ok���aR�!�`�(i3�S��Y\&U�)j�S�mJ�0�6�!�`�(i3�tU,�Ql�	^���y ��-O$U1tSjv�!�`�(i3�(R\֎u��w�`L�h��=��޵g!�%=F�=!�`�(i3^	QW�Q!r�{F��#��g�+C��s�t}�F��<�����xb�ݚ�Н���F���K�&�a�M����*��q9+t�}�ݚ�Н���F��=�?��3�M����*�'�^�����ݚ�Н���w�w:�!�`�(i3^	QW�Q!r�{F��#��g�+C��sJ�A7���ݚ�Н���F��=�?��3�M����*��q9+t�}�ݚ�Н��H�����\�2��s���1�, �y�`��vN*���k� ��$J�L�l:�
d�rP&��dGL�F�z�>�/�O8���6�d`̮�ӋH�RtV�^!�`�(i3�b��+N���ˇF}<P_�H�RtV�^!�`�(i3�%t̓�@���{
B֗M-k��%)z�
3Me!�`�(i3��w�w:�!�`�(i3!�`�(i3�$�������_j���=n��c��>������!�`�(i3���F��O��ݚ�Н���'T���+�%�эȈ]Z�����q9+t�}�ݚ�Н��Ra])n#���{�@��$J�L�l:�
d���:����j�V��veK�	�$V�#o�]�ʄ����n�0R��#���n�zq�����X� 2!�`�(i39�6M��",oMG~�>y�pA��w��+-��, ��A�Y�
���3ʩm[s����������)e��e���N�ScG�\̒=��!�`�(i3ݑ���&�d��ҟw���Z9�+	�I�e���U���}Dq�f�!�`�(i3�\�2��s�pRF�E����{�j+�j)����r^!�`�(i3T#�3�["�7#1=��*�Ь3Ǽ��״$(�>g�!�`�(i3��F���K�&�a�M����*��q9+t�}�ݚ�Н��Ra])n#���r����!�`�(i3�$�������_j���H^�h���i��}Dq�f�!�`�(i3�\�2��s������x~>#�+#��]��}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4���ݚ�Н�����,����'	�!�`�(i3�\�2��s������x~>�"ª���ž_�F��H�����J�g�*�7�~�k�_�mS8<�n�ݚ�Н�ݑ���&�d��ҟw���Z9�+	����3��[<�m��I�!�`�(i3�\�2��s�pRF�E����4�'��'�Ƀ�?PA������B!�`�(i3x�j؀O��(�\G�@�L^�?����NM���
�:qEp'{w#/ B!�`�(i3���{�@��$J�L�l:�
d���:����j�V��veK�	�$V�#o�]�ʄ����n�0R��#���n�zq�����X� 2!�`�(i39�6M��",oMG~�>y�pA��w��+-��, ��A�Y�
���3ʩm[s����������)e��e���N�ScG�\̒=��!�`�(i3ݑ���&�d��ҟw���Z9�+	�I�e���U���}Dq�f�!�`�(i3�\�2��s�pRF�E����{�j+�j)����r^!�`�(i3T#�3�["�7#1=��*�Ь3Ǽ��״$(�>g�!�`�(i3��w�w:�!�`�(i3��l�^!Fڸ�>P��=����h��A~����>������!�`�(i3x�j؀O��u�>����Cw�Hm��!�>!��!�`�(i3^	QW�Q!r�\1^O� �Xz���%��v��!�`�(i3HN��R��bP�63Z�t���%>�rGO�D mWN!�`�(i3�ݚ�Н�t�cz�C�55f�)�}!�`�(i3�tU,�Ql�	^���y ��-O$U1tSjv�!�`�(i3�(R\֎u��w�`L�h��=��޵g!�%=F�=!�`�(i3^	QW�Q!r�{F��#��g�+C��s�t}�F��<�����xb�ݚ�Н���F���K�&�a�M����*��q9+t�}�ݚ�Н���F��=�?��3�M����*�'�^�����ݚ�Н���w�w:�!�`�(i3^	QW�Q!r�{F��#��g�+C��sJ�A7���ݚ�Н��H�����\�2��s���1�, �y�`��vN۶&��L�H�xѴ�� ��0>!XM�#�yP��C��?�T'����M?��y�!�`�(i3��l�^!Fڸ�>P��=����h�5���`�!�`�(i3�_��>νrj�V��v��=����n��뾦�!�`�(i3�_��>νrj�V��vG�?-�D%��v��!�`�(i3�߆�p�hع��)/^��>&S�XQ�u�j�fKÀ�:����j�V��v�Gj7�uz_�mS8<�n�ݚ�Н���+�t2�4��A妡��M/*�3҇	��*��O`�� \)!�`�(i3x�j؀O��%c5#	�.� ����7����|e"!�`�(i3x�j؀O��(�\G�@�L ����7����|e"
�:qEp'{w#/ B!�`�(i3�%t̓�@���{
Biۧ˺�s ����:N!�`�(i3T#�3�["���'(��Cw�Hm��/��kOT!�`�(i3T#�3�["�7#1=��*Cw�Hm�̊��NM���!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �m�ڨ�hծ�ݓ�W���=�����]s���D*j��'T���+�%�эȈ]Z�����q9+t�}�ݚ�Н�T#�3�["�7#1=��*Cw�Hm��/��kOT����l��-4fV���d�ވQ�:�G��Hb� h�ҩι�+�t2�4��A妡��M/*�3���X�zK;��t��:!�`�(i3��+g^l��~��w3*)/�k�2�i�:`�+Py�b�G2!�`�(i3��jVѭ@!�`�(i3�%t̓�@���{
Be���C�������y�!�`�(i3^	QW�Q!r�{F��#��g�+C��sJ�A7���ݚ�Н�$f��_Ub�F�S�1 �(*�O�qe��0�U���>e���̰�!��U`�PW}D��ɍ��Wsp[��X��=@'ѥ���F���K�&�a�M����*��q9+t�}�ݚ�Н�T#�3�["�7#1=��*�Ь3Ǽ��״$(�>g�!�`�(i3x�j؀O��u�>����Cw�Hm����x�a�t!�`�(i3�;b�-�2��Q������}�	76�&�φ��<�6��(R\֎u뽀�%���eZ?�[�-q�\E��09mh��n���K׵��φ��<�6�@a� ����C�'�ąC>��Ӛ��S�J\7r��*�t�>��G���\���F�`y������T�8k��.ͥ�H�RtV�^Q� �_tt��`���`E�g�������(ӈ���m�r����̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l��|<��r�*���u��
�a��o���H�RtV�^q�\E��09mh��nFe��1��'��L�㜯}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M�c�r%�7�i"T��]���'z��F�c�r%���_��J���J��ۍb�o��_�Rv�䩲$����#��i����+�^n=\f�5>�OS�3M��e`�!��:�r$ɓǉ�.y�U=������&G�wӨj]h�u�#�$IX�E'���dN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H����|��sQ�G����)�
�M?��y�!�`�(i3Q� �_tt��`���`(C�d)խ$�����z��ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;�끓��~�Lu�#�$IX�0w�Ʉ����'z��F�c�r%��Y��a��G�}��ɣ ,��rQ��NۥUn�`��c,�Zb��8��Ս��Z�å���jVѭ@!�`�(i3!�`�(i3!�`�(i3?V��j�c<o�;)�y�Pt��`������,�ǰ�,l�=�;+i8�
B�*�x�uD�b�Y�c��r���i3a��o��_�Rv�䩲$����E)e|A��`���φ��<�6��7�癆cgR������������ h�ҩ��(R\֎u��Y������y¹߆�p�hؽ!�M��9�a>*<UB3 �~k�%�������&Gݑ���&�dw�c��l�,�ĉ�Iऱ�ҟw��Aɠ�T�nGHN��R��*9x���С$�)�vx$�Qo'2.�t�|�AS�댿d���;U�a�(���Ņ�F'φ��<�6�@a� ����C�'�ąd�G}%����3f��gmJ/���'ž1�|��P�:k& ��-����^	QW�Q!r�#✲�@�G�-�6�T�my$�N��o�/���;�̢k���"��w6�0��ɗ��zi#Y)M���Fe��-����u?�:�H���z��l ��8��GM��-�����_��>νrj�V��vJ�
�M��}��u@:b����d�	��uc���F��O�}�	76�&�� Ӗ�t$�)�vx܇1~�}������P}Ѷڶu�7��9;��ˉW��	]�	�U��)���Y;e�iK-pm!9�>��n4s1��7�癆cgR������������ h�ҩ�x�j؀O��w���B}�#QSU:�����|e"\���>����!�|Dk���������|e"\���>��XKH��Κk���������|e"O�.����B<�L�V_�I����~u/��kOT��$���͜P_�_S:g�RMm�o��'����u��r�助+g^l�>&S�XQ�2-�#?C��%�э���T3�!�W���b�0�Р�(�V��M��:�j?������e�����=;
����cp6Dq���e������L�$�K�dߧ.�go� �e�d��rp"n���m�z��P��4AL���c����L�{v{��lw	U�d�#�b0�:�#�k(��Ě���aT��3G4��������d'��",oMG~�4��g%j�V��v
���=bk�Bӫ}}5'G�+R���o��_�Rv�䩲$����E)e|A�յ[+8��r$ɓǉ�.y�U=������&G��F���K�&�a�W�^�|��/��kOT��$���͜P_�_S:g�RMm�o��'����u��r�助+g^l���b��M�4��'���K�&�a��(u�A�HN��R���ء�I��߸��S�ȌA�GIp�7�,��n6�o8:4�I���c�90Mj�dL���èVxjzӝ���w3��׍�&�U��f��_��>νrj�V��v�k�n�=���b+}y[�k��^�1Aj��t�35L��$
8��2�ֈe1tSjv�T#�3�["�7#1=��*���3n�v�j�V��v�Ȯ�F��}�	76�&�� Ӗ�t$�)�vxƮ���i�f�%�эȿ�O|����\�2��s��t��������d'��7#1=��*?�4V�I�\1^O� �n}沁,yO�a���R9��φ��<�6�@a� ����C�'�ąd=��¾ȼ\���F�`y������T�8k��.ͥ�H�RtV�^�\�2��s�RdE�̈́|J�A7�伩���@|��璓�c�������t �[l;M?��yЮ_��>νrj�V��v�.R�x�j؀O��u�>�������W���Ě���aT��3G4����~��cǞg61 ��.��Ã���HXy�<ry��!����T�[��.��Vr���J��:�����#}�{�\ٿ�6�P]M\I��A$�P��O�@י����z��q�`���φ��<�6��#}�{�\ٿ�6�P q��j�J^�'ž1�|��P�:k& ��-�����_��>νrj�V��v�f0� ���nF���<�W�.�P�	��
�Q�}�k��^�1Aj��t�35L��$
8��2�ֈe1tSjv��H����|��sQ�G�Yu�������&G!�`�(i3x�j؀O��{dOCe�@)X��ėd�'��L������*C?7)D�[
�:qEp�;�P�t�5fĉ>99��A0ok�׹�>�)� H]o���B�m��d�uu�w�R���y���Aw9��x�S�ӄz4��+n'��hE�8�Vg��L�*�!��ҷBcB8��I�G�p�P4&Ƒ:2�c<�^<�H�W+��W��\�2��s�ώ ���]q�;&=7�kJb�z'hۉ)��d�7�qĜ���,�ǰTm�v��G�kv޶Glݓ#���照�'�u����Ƶ�ӫIX0F�MV�ҁGG�K�BN
\����+�^n=\f�5>�OS�3M��y��>>�����qD��=a�^7�1tSjv�EOJ�uxm�	�����e��0�U+�qbp@��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#;�j�����g���Qrf_�mS8<�n�ݚ�Н����'�u���i�Wg��+Ut������F��O�}�	76�&�� Ӗ�t$�)�vxV�/e�,�5���)D�ʵ�b����:W�����t�T��?E-h���U���e��_	�Ƽ��S�J\7r��*�t�>��G���xjzӝ���w3��׍�&�U��f��2��}����+�?nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r���_��*��jC��6�g���7t��'�1tSjv�?V��j�c�4���<t��&�*楉��%>�rGO�D mWN��Ě���aT��3G�IX0F�M�}��u@:�K���w����s�`夊�V�%�1Bd�.e�R�;o�� ���nF��kJ2�,����Iwl53�e�'{w#/ B!�`�(i3!�`�(i3EOJ�uxm�Pt��`���,��7-oc����H�}��ɣC��r�"���X���&R`��c,�Zb��8��Ս���3�vd'{w#/ B!�`�(i3!�`�(i3!�`�(i3\���>��XKH��ΚM��%�p@!�`�(i3�mJ�0�6��A���A3�p��(�l��c����)e��H�d٦�[*�,��7-Ə����|��&g",oMG~�j�ā��u}��ycĢ�<�..�4����Y<�!U���t�T�@$ �O=� �e�d�����`��u �e�d�������x����0��G	I���e�!�`�(i3!�`�(i3!�`�(i3!�`�(i3��f�,�k]Swx�x�K_��:��8��yP��C��?����FCA����.���<�ry^�!�`�(i3!�`�(i3!�`�(i3��l�^!",oMG~���	o%����(R\֎u���j�p��ݚ�Н�!�`�(i3!�`�(i3!�`�(i3���̰�!�Xy|�W�]��(j��_~s�8���v��ޫ��w-��n4s1�%��W���ff2��O�ܬ!'B�}<���E��D�G�&ց�*�8a�qK�X!�`�(i3!�`�(i3<�6�Q=�-��	q[^�Ր�rj2�ݚ�Н��(R\֎u�=7�7K�P�"ª�����}Dq�f���M2�M�;Ss]�k������8#һ���}�}D��N�W{��ǖN┛Z��p�7�}�!��i|�rBY�",oMG~�Յ$�O&�#o�]�ʄ�< �SS@�
�رjwc�';��#j�ݚ�Н�EOJ�uxm�}�Z��y�&TL�b��!�`�(i36S� �*���8�� ��V���ޕe`�!��:��w�w:�!�`�(i3��M2χ����a�)P<�ܓ�Y
�:qEp�;�P�t�5�wӨj]h���z��l 2�����4ƍ2���lČYw����~q�_e��!�`�(i3!�`�(i3�e]�#�?5���n2���}Z�
d~�r:]���!�`�(i3oв%u�K�>&S�XQ�Q��rj�_\q:��gT�-�c�I�gV!�`�(i3�%t̓�@��܋�n焞 ����7�[���n<�!�`�(i3�B�],Z(i���Fz���l�^!ЙMǿI?��6�a���}��Xׇӭ��fĉ>99��A0ok��ݑ���&�d�����l9�̪=���z_n�ԁ%m�\�u�K���/Sg�Dzy���(DY&���;�jmT�#�G�2ޟ'H�\�{\�n	ͷg�?������2|Q�-l�;�CJ?К�-����!�`�(i3|��sQ�G����7E�׵��vH<�6�Q=��[K�9MY�^�9�Δ
w!�`�(i31���~�wӨj]h���z��l �"�Mg�ƍ2���l�HN��R��bP�63Z�tq�\E��0ÿ����Ԗ&TL�b��hO���2��bY�[�&O_\R'�I���gT!�����p!!v*!��r��  �wӨj]h���z��l 2�����4ƍ2���lČYw����[�ǥ<^y!�`�(i3!�`�(i3�e]�#�?5���n2����k	�����l������l����)/^�蜬�^���'ƃ�3�Y1tSjv��wӨj]h���z��l .+�N�R����|e"��w�w:�!�`�(i3��M2ϼI�)�ݳ���b+}y[���%>�rGO�D mWN;�jmT�#�(R\֎u�,��7-� �9�!�Q��s�s�{��ҽ��d9=���u��r���2��}�����U��f���0z8#һ����~���U���O@���zxC5�h3]�< :�!�`�(i3D"ۡ�
",oMG~�>y�pA����v[v%��%�э��XW�G�<a��o���H�RtV�^��l�^!ЙMǿI?��6�a��)P<�ܓ�Y!�`�(i3��jVѭ@!�`�(i3�%t̓�@��܋�n焞X��ͷ(�-���|e"fĉ>99��A0ok�Ra])n#���r����q�\E��0�p[nۈ�I����~u/��kOT��+�t2��iK�D�b=G�6�!~�%��v��!�`�(i3�5ߧE4��!�`�(i3|��sQ�G���I:)�/��kOT(*�O�q̑`�_!�`�(i3!�`�(i3��I���x9[���[�� �<4��Kƾ�*��Aڬ&W��%�э��XW�G�<a��o���H�RtV�^�u{*�C<��e�����(�G�$�)�a��o���eo<����UEv����UrO
���,|F��w�[�?Ve�|9����l����x������Z��������&G!�`�(i33�[ד�������l9�̪=���"��ӌ�r!�`�(i3I�c��C�p[nۈ�q9+t�}�ݚ�Н��wӨj]h���z��l 2�����4ƍ2���l�.Y΄�l�j1���~!�`�(i3(@X~�H:����dܟz�-��h��ƍ2���l�!�`�(i3��M2�}'p5���s)P<�ܓ�Y!�`�(i3�H����fD��j��ه,��7-� �9�!�Q��s�s�{��ҽې���xQ�1tSjv�!�`�(i3?V��j�cC��6�g��3�J��~m��}Dq�f�!�`�(i31���~!�`�(i3?V��j�cC��6�g��3��	cA霯}Dq�f�!�`�(i3�5ߧE4��!�`�(i3HN��R��bP�63Z�t!�`�(i3�ݚ�Н��5i^�����d��&�A�k�������!�`�(i3���̰�!�Xy|�WCw�Hm��/��kOT!�`�(i3;�j���������^��b+}y[!�`�(i3͒t�]��/",oMG~�Յ$�O&�#o�]�ʄ�< �SS@�
�رjwcgWaU �IH�RtV�^!�`�(i3|��sQ�G����7E����NM���!�`�(i3��jVѭ@!�`�(i3q�\E��0�p[nۈ�q9+t�}�ݚ�Н�fĉ>99��A0ok��
�:qEp�;�P�t�5!�`�(i3;�j�����ۥ�Y�m���NM����Ra])n#���r�������̰�!�Xy|�WCw�Hm�̊��NM�������l��}��>�u��M��:�j�7t��'��uΜ�6Ä!�`�(i3��M2�}'p5���s)P<�ܓ�Y!�`�(i3��jVѭ@!�`�(i3��;��L�ז�1�, �g�f�p~(ŐV(MH��C��|���8!�|!��[��-����!�`�(i3��M2�}'p5���s״$(�>g�!�`�(i3��jVѭ@!�`�(i3��M2�}'p5���s)P<�ܓ�Y!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �?V��j�cC��6�g����$�\%e��}Dq�f�q�\E��0�p[nۈ�q9+t�}�ݚ�Н����F��O�/�"����V(pyL0DMlE'�! ��l�^!ЙMǿI?��6�a��)P<�ܓ�Y�wӨj]h���z��l >c��?�%��v��!�`�(i3|��sQ�GD��P��Z�q9+t�}�ݚ�Н�;�j���Ѐ�K����$�\%e�E�i�m}6�4���n��Fr��j�p���"�|��c��@��Y?;t|��JL�����d�ШM�EfS�	Q���f����.����{ɖ!H�mIZ�q��6�^��ݗƩ��F�z��b�m��HNf��q����Н�:���M��:�j����j&G�p�pU��mx�j؀O��)����bXem5��3'!�`�(i3!�`�(i3���D4FF^�i�H��,����I�S&��p;�E,	P�QUH6"�w��B�j���;�����cl���,��7-�B�9��-4�@	�u�a��4	_��%�э��XW�G�<v"��1^�!�`�(i3{�d"����	�,�2ZL�ԸK�F�W��	]�	�U��)���Y;e�iK-pm!9�>��n4s1��7�癆cgR������������ h�ҩ�&����(Au.$���k������8���[{/;tiND�S���/9�=eSe.��a��o���H�RtV�^���{�@|�;�Ojz�$�AՁ�Va�ir�\�2��s���z������r��$��0�'z��h{���kS&Q��gVdxQ,�,��7-�B�9��-�Va�ir�\�2��s���1�, �~ܙ<�Sd��Pt,Y�-�_{sxJ�a$�Y ��M�
QC7�T���Ek���,���Ě����E�i�m}6O�D mWN��ܐ�}Ğd��5��4PB����A#��Eo�3�IX0F�MV�ҁGG�K�BN
\����8-|�D���"sS<GYqcHTX�';��#jx��7�֕iK�D�b=��L4�����Ǉ�y��}Dq�f���_~s�8�c�kg��k������8���[{/;tiND�S���/9�=eSe.��a��o���H�RtV�^�K�&�a������kO�h|O��ЙMǿI?!����a�};�jmT�#�(R\֎u�{��b�b�*#o�]�ʄǑ�+�/Z }�Z��y�w���;�j����" �,G?�x{^4��*m!�`�(i3��_~s�8�c�1���7�?D�8���k��^�1�K�&�a�/�dI{�8k��.ͥ�H�RtV�^���#Ge<%��a����z_n�ԁ!�`�(i3�֊���}�Xy|�Wcz������Ě����E�i�m}6O�D mWN��ܐ�}Ğd��5��4�iK�D�b=C��CFv$����Wj4�RtZ
Xgp�(R\֎u�=7�7K�P}��J�0_�iK�D�b=\#�!V5ȑ�(R\֎u�=7�7K�P�Bv����`��)e��[�<� <��^���H> ��+�O�XÁ�p[nۈ�d��-��!M�2*详p*�з=I�^$D����(R\֎u�{��b�b�*}2��L� q��j�J^!�`�(i3!�`�(i3myC�0kc��g���Qrf�Va�ir��_~s�8� ���3�<<��lpЙMǿI?��g�F��6�>Jj:&ֲ!�`�(i3!�`�(i3���[�Q����U4����#=�Q��s�s�{��ҽ�1F#�֞q��KVט$����dܟz�L�[\�"��jVѭ@!�`�(i3!�`�(i3����(��e
� <"w���U���LQ�/8��u��m�byBH�}�x&���Z�߲��-��F�M��:�j�r�~t���َm(5!�`�(i3!�`�(i3!�`�(i3��yb�	�����u��
�b~*��s�!*Ĭ����x��w����iK�D�b=`u0�F��a�D狹�����zԏ�E��e�����U|�W�˷�I���!�`�(i3!�`�(i3!�`�(i3�%t̓�@���{
BfxQ�-V�N|~�.�u���r����!�`�(i3!�`�(i3�,��7-p ?7�7�"Р�(�V��M��:�j�J�a�sb ڥ����ȾmyC�0kc���Ø��4��Va�ir��_~s�8	0X��f*��<<��lpЙMǿI?��g�F��6JJ ��iG!�`�(i3!�`�(i3�F���ᘮz��l Ю��U������2|Q�-l�;��5��t�;��Cٯu�Xy|�W�����z��s)l໶�,!�`�(i3!�`�(i3kǿ�E�Q�C��6�g���7t��'����+���b�6��R��J����;4�zu%��0q�#�<���H��K49;��Cٯu�Xy|�W�4Adq@z!�`�(i3!�`�(i3���D4FFo����>�/|��sQ�G�Yu���km�������.���n��Zn���EU.�Bft>��#o�]�ʄ�< �SS@�
�رjwc�Va�ir�K�&�a�/�dI{��8������k$ !�`�(i3!�`�(i3Р�(�V��M��:�jE5�����]����0��G�|G�N.�N�ܮ2�k���98ޥ�j�V��veK�	�$V�#o�]�ʄ�	]�k��,���^���'ƃ�3�YЄCwc���)e��e���N�Sc	z�{�eM���8��Ս��%�r� �7���U�� �e�d��C=2��km�������.���.����2�hY�%Ͻ���U`�PW}��[��o}L��@�.�'{w#/ B!�`�(i3!�`�(i3��ɑ��Gj�Q*��a�,��7-P�OrY4�b~*��s�02�ok�+�g��{�峉%�2��)e����U����+�Va�ir�X%�;���s��v�c�e9�h2B��͵h.��r@�A�A
i�eL!�`�(i3!�`�(i3!�`�(i3x�j؀O��w���B};���{!Ae0�@\}p