��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G0��@h ���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω������?9X�1�Z�U���T��ײ2��>���^k�/7�?1�(�c��ly[�$D֍C95^T��6\Xa��7��Į�N��=i�@x_\q[�@�0�I���j{�N<��;��� B]�pE���	x]̃Dj#^Da����M���v��W�&��v�=�z����)�,�˛D��w���旴4�����<��a��rl�ʩ{�Bfळ��)���X�$� ���jǎX������n�q��}�p� �Ñ�]�*�p�㈍x�!����Y�f��a�Z��Vb$���N[E�=����tL��	Z�G�a}CK�fC���4�O�"�F�È���_�O��<$e|����w'��1�:�Ω������?9X�1�Z�U���T�����\�4�sP	�b\qB��������"^Y怄����v�~�MUs a"�x���2@�+���c�#s�0���!Z:���:r�a�u�����!�M��E����F
r:�����u��w)�S�5� �7��Mv�9*���f��^(��f�)y�8�:r&@��=��$얃�rb2 �Q[1I�����w'�\�Q�3M���e�t��yn�	� �x�m��n~�q({L�51��;����'��%Ճ�86���H�aF��6��I���j�r�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�E�s��bc�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�y���}�ZC��aNvA�;��>Oʉ�~09h�i�k1i�f1?�e�Bw�M�?_W�\I���A#|��[�m���w��L�����'�{b�2"���Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ��4Z��ʬ�,I\�Z˻r���V�>!�/�7��u���nEA���e�q�L�Xڈ*-}|��ι%9��oGo�Z�J��ݪ��4Z��ʬ���Ӿ���	���q��q�©�����<��������/�����,��B	hI�ˋ��b�ӝ5�T�@���k�փ��㛋��X���`��.�̀�I7��-5?�1J&�|D�e�!���QI�D/����ʊv.s/�B{�o
�Y-�E�f�}�=Ll�����,۽���}i�@�5�}�]���x�]�V��7��_��T��!e����\G�Y�)��Y櫧�7*9uu"�,�>E��<��z��}�0z�cUL�n����4���á�~O�"j���b7|#9���[�t��#���j;9ekN�By3��<Z鎬�������(���P����ˮ��lC��U�T�\ ��+�_0c �Q�P��
S��j���0z�cULjaGkƊ~F˯�+)�"j���b7|#9���{k�h�+�����
L'���Xw�j�7��ct�:��RE��W��_�ړ8���/�z&v��\��t������S�)37J*u>����C�/����o<��z��}�\w��0]Y��
�iC�o��C!T*�q���U�ЂDa��(O�J,���Z鎬����F�71�B��O1��m<S�)37J*u�񁫴}2��:��ӰӒ1�:�Ω�>�����V5�"Bb]1]M�Kz,M� ?ҡ���y�E�nwE��S��}|��XH�����,>$+W��� j�(����5���ռ�j��I���j{�L�Y�͋�<q��?!y�A��-|�t��-?dȵ�ixUS�/��A��갖��fb��иܖ��5�rP�'b&ʝi3��,�&� +J�����|����OxtX+�Yo��Ⓖ���á�~O����}���7�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e,%�0g�������DzL��L96�`6�CY���<�I����"�*�şxˏ1"Ohƪڈm�d�٣��c�A�L'R�o�����5�%]���a(􆿳���2����.〧I���2��� �� Ϳ�$��0z�cUL�n����4���á�~O�"j���b7|#9���b!��u�G��ô��~ ��ç�Y�{'%s��.|Z���I7��-5��6��	���`y����@����gGWm?"<����;F5@0�Z鎬�������(���`$�P.eE���lC��U�T�\ ��`��K Y���S��I���;E�@
�����8�l��m�f�$|�/|�z��#G���q����<�6�Q=s�׾8��Ρ�Q��nT��Q#>[�/+mQet!�`�(i3"�,�>E��ʆ�In��tT?�7G|`~�Y���(�}�Π�cC!�`�(i3�i3<�f�D���X���`>���������Y�l,r\����"�,�>E��ʆ�In��t�_�R�G�������b�Xϋ?@)�ak�m6=]A��O�T=�4e=��-��Y
���t�9�,��Zt%��m&<Z�#�j���0�5tU���+�J��U<o^.K�}/��<Ӭ�hDJ��3Y� 2��4�b��{�P}�зq8�Ј)w�<�_N`E�cvR+��}Dq�f��d �S|�b��{�P}��E����F���8�TP��@E�`�8���&�r��SQQ���bK�&М��!æ�4];ˍH����TI��Ԫ,щ�">k0��Wp7�:�!�`�(i3x�]�V���t�����[F�a�+#�n�%�<�'`ٲ�)�ak�m6�a�\����8x<�A!��=����t��cg3/F�C����Eb@2*��N)w�<�_NX�ʟ�3���M&������h�? "a��Q�V!�(�x�]�V���t���	h�Tn��<�6�Q=>V�A�$��Q��nT��Q#>[�#�@�o0!�`�(i3!�`�(i3�i3<�f�D���X���`>����������o��,�Xʚ@h!�`�(i3�i3<�f�D���X���`>���������Y�l,�x�6�
X!�`�(i3�i3<�f�D���X���`����"�I��j&���.���7b!�`�(i3=]A��O�T=�4e=��-"w߻Y��}Dq�f��v1a{J�^�|n�M�!�`�(i3���D	��U�l>o��|���JLm|�hDJ��3��`%��nx{<qH�~�!�`�(i37�ܥ��2�A�Jr���CVF��g�M��p���!s�;�����,�Xʚ@h�E����F���8�TP��@E�`�8���&�I��j&����bK�&�B�r��=]A��O�T=�4e=��-Y�VN�=�ԃt����}�b�Xϋ?@,�Xʚ@h!�`�(i3x�]�V���M�K�=g�H{g�q� �zbw��(����~w?)���0�g��^�}#4];ˍH��\B�����g�q~[{Q�Q�.�`��S�ƥ���!�B�r���E����F���8�TPm=_g}b��t��ީ�%�Ӫ�p�B�E�!�`�(i3зq8�Ј)w�<�_N`E�cvR+��}Dq�f���R����a�=L!�`�(i3���D	��U�l>o��|���bǬ�=SƏw0���wN��0]�k˗S�d�"�,�>E��4];ˍH����TI��Ԫ,щ�">k0�ު�p�B�E�!�`�(i3���+�J��U<o^.K�}/��<Ӭ�/�"�����_G��?'���o��!�`�(i3�a�\����8x<�A!��=����t��cg3/F�C����:�,x�~7�ܥ��2�`e7��9���I^Ɍ؝�hy�/B/���^!l���Z1�:�,x�~x�]�V���t���CՐ3��F<�q7�0������v�e����~D̤"�,�>E��4];ˍH���*�Yb}?iRPsNR�r�_�L���+�]�iJ��@x��D���j�C�6̓126��G}!�`�(i3!�`�(i3x�]�V��h*w�N��M5�v���Lꂐn��/�Ζ�{Q���TI#!�`�(i3!�`�(i3!�`�(i3�a�\����_~�7�(�6k�4d����1�so��d�a���A��`�c1+��H,�^��'�l>o��|���&l@��,щ�"1��tζ����u*Q�!�`�(i3!�`�(i3зq8�Ј)w�<�_N���i�ꜯ}Dq�f�p 26af<�B��+ H!�`�(i3!�`�(i3=]A��O�T=�4e=��-j0��.@.��}Dq�f�p 26af<56ND���8!�`�(i3!�`�(i3=]A��O�T=�4e=��-j0��.@.��}Dq�f���CZ���%gɚ��Ol2!�`�(i3!�`�(i3�i3<�f�D���X���`����"��L�K��%<7�`+Al��R��!�`�(i3���+�J��U<o^.K�}������9b$ɠ����T55�\H{�U0X��~&����}Y{!�`�(i3зq8�Ј)w�<�_N�ҕ�:9)5?iRPs�;�.A�ى�P�p ��=���=���a��z>�n�SS7�8�8�&�3Z�K�x�]�V��L3yJT�`&N�V��<���O�;:�<����E��~@�k��ϳN'��+q�3[�u8���/P?�c��t��L̿��$|�/|�z}��Hn�[�57�0q�7Ê7�E�4'���Xw!�`�(i3!�`�(i3!�`�(i3!�`�(i3)��� ��1���J�aK�#���o)��B�ӮY�E��vNd�)ir���j:N�By3��<Z鎬����a�gN�3c!�`�(i3!�`�(i3!�`�(i3�����C�#�ҒIs{m�А�V?������m���B�Nopa�ǂK[���#<��z��}�z�-~BLI�!�`�(i3!�`�(i3!�`�(i3V����(n�	u�!��qő��{��1݁mP2<WV��
i�c�r����P��7Ê7�E�4'���Xw�j�7���1�)�c��,0=]^	�&�e A7YzE�ˇ�h����2�[Q	��
�Q�}#�ҒIs{Y��~���B�No?V��j�c�m�LT���<��z��}�0z�cUL��լ[po��vf���g��U-�eq����9�K7͍��ճ��)�ȓM�Me���섫�So#�[�}��|SM0.�J�a3mPykIt���	�]�!��	Ǹ�y85�&�;���
j�T�ܪ;�T�\ ���:5A��p��1����lovMVgd�a�"�
�������iA'R�	�o��C!T*Y�{'%s��F���kU0F�o^�V]��}��ł�!r�dN�<@Iv�,.9������:5A��p��1���#Dfc[�gd�a�"�
VA�ڦ�c4G��.��e��n00�8��P6�Y��\���(����A-u��6�0;��ȓM�Me����ΜtȓM�Me��x�2�Hxl�� ޘ_�9��\�'�������>Q��?qr�)�b!F��>z�����&�զ2p�$�W��	]�	���F���X:���m����x�s��J���Ş|H��S��q<� �77AƐ^�87��I+�T���B�H��y�&؏R!׻�p���f
�@"��wҦ�kQW֑��bk<����-I���z�S��Ԥ�ء�wrq��c�\VȓM�Me���T��G���X��4tΘIy�����OyQ���؟�-�X��_��n��&�PRn%�bM��pK���|�"u��,�ttT��4��G{Z鎬����=���ޒC>��}Dq�f�d´NA�*Z<��z��}�<ͧ�:|zG�_h��� л�?� �٠FӮY�E�/�^; �
�0S&",f�e�0�؍�3Ϟ��M�+,[�� л�n&����_!�`�(i3!�`�(i3���y��lD�U&"���+c��k��Vj����C$��*V�ֆ�˳k�L��<�6�Q=� 䉇o�M�· ���4!�`�(i3!�`�(i3	g u�XI��ׅk��+ņ\.���(b�rq��c�\V��=����t�6+W�آ�{l�f|��:2QYeƈ״$(�>g�Y��j3�����o�g��ҋX����L$�����/���%��Y�i`YS������I��q���Um��#��*y��+�^@��#	Ͼ7�Z#^L�)�4)	���E7��I+��v��q��y�&؏R!׻�p���f
�@"tL�^VG��T_�[�S{\bE����25��X�N̘Ľ|�	���c�.D٣��&�զ2p�$�W��	]�	���F��qJ�?�̃�*�`��n�E�T����X�=���P�;�ȓM�Me���섫�So#ȓM�Me��x�2�Hxl�� ޘ_�9��\�'贅���Ǯ0��]㯟B./�<ĩku��j�,�J�2�|bQ��� Ǐ˨�g����K���=
��P��bE˧�<vr0�����i�é�I���z�S�*��iMOP;�
2�P�nlH�Ir�VU������ڑ�eo�]�!���\B��V���|e"{�7��4<��z��}�<ͧ�:|�>d�g�KSƏw0���:ʽ�f��x�	-���]�!���\B��V���|e"�'�al��p���K酦��{l�f|��:2QYeƈ�	�����Ζ�{Q�]~'�H��{l�f|��rs�i�Vw�C�-�]|If">���%�o)��^�V]��}��ł�!r�dN�<@Iv�,.9������:5A��p��1���z\�=d�#Q�
_�J�g�J�LQ��w֚S��~G�݈,��S�)37J*uc�A�L'�i����
��8�����x��3�a(􆿳�tP"7��%e��0�U�S{����<�6�Q=�qő��{�q��7-]P2<WV���Q�pA��i�����R_"@�v�{�&7��U-����`kv#`ʽ�V	=�7G#+�Ǘ0z�cUL��լ[po��'N�*	�g��U-�e6R��h��MH��WZ�mN�2߄�84 �Y%��(�
t��Y�{'%s��F���b��8��7�v�ԯ�>cg�`��섫�So#����hѓ؏��ǖ�!<��}�u嶅 VU+I���!�g�%���ۂ�3�����U�8"�,�>E��Rݛ��%�5��lW0۳�*ȑs;��|B����k2��� �����!�`�(i3!�`�(i3!�`�(i3^�R���c+��;�����$�`V1��eX�:&���!�`�(i3!�`�(i3!�`�(i3!�`�(i3�gKh�ߕ�ő̓Vo�ArV�b���0��!�`�(i3!�`�(i3!�`�(i3�I����~uոA2t\�����F9�@�8
�O��Gs�m�6�o8:4ڎ�\��q����+�^n=\f�5>���j����v�۲=�k2;�jmT�#"��w6�0��ɗ��zi#Y)M���Fe��-�����2��}�������K!�`�(i3!�`�(i3!�`�(i3J�a$�Y ���q�}�:�yB�x�$f��_Ub��7��G_��$�)�vx��j����8
�O�h=<*��q\$�ҞC���!�`�(i3λF��|�o��_�Rz���n H��èV#�աl�P_�_S:g�RMm�o��'����u��r��q�\E��0��)(��8�!�`�(i3!�`�(i3!�`�(i3�I����~u�L�s;SF`L��n��p��b�Bϱ��5?�&P-��:���Y!�`�(i3"<�GU8o_�mS8<�n�ݚ�Н��tSk�N����C.�u`oPϞX�o|3��b�Bϱ����m�#Y�N��b��?)ݝOv%:�yB�x�fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vxo���.��@K&��H6j�"Hs��.�X�Q�H���sd%4Ӥ�鏄�!�^�����L��>���	��=�w������K���'OWb��]��F�,�֏��9�GͿKR�7h�,b0V�u�Q�ݚ�Н����2wG!�S�@�]_LO���׻�t�"hzf�?ǉ�=�+�H>�?ۭ�����b6�ŏ ���N���B
���?�Ho2��2�n���mv��6��fC��T�z���,}l#�>b�eIG��Q�q>x��b� OEfVNNaJ �!,¥�����Ј��wf-��w¹��<d�,��L���D:���̒!٤���!�`�(i3�F�7��Y�
�cc�V��ݚ�Н�I:�K�R����4�txj����R��á�~O��&�C�/:��+���<eκ3*Y�AQ�0G�F�r�f�t�Jb�[���B����n��e����kn4@Q�/�!�`�(i3����@�&8�,������	�;�ݚ�Н��'�al��p)�ak�m6�0��"��S8��4�J	~�ւ�J䏊Zt%��m&<�,0 �����X;p`�Z鎬�������(���G�n봈2=B7Ԅ���s�٩�����w0�H��bf�?ǉ�=���K�Ȃ�H��bf�?ǉ�=��9K��r|�����KM몴PBoT�ݚ�Н�� 䉇o�M�x��f�?ǉ�=��TBd��p!�`�(i3�d�)bU/�'5�����@�_&!�`�(i3��%ў׫��8q�/�\4L$ֵ�)�ak�m6�e�-3��ݚ�Н�|�� Cy�6j�"Hs�Cx�V����c�RjVU�簦D�L�x8�̹�y3����&=)X���37�˱�5�ݚ�Н�{�"���ڥ9��[;�h˒�Ӆ��uՇ�OD� �B�S|�P�DM몴PBoTη��~�������
L'���Xw�j�7������}0`a(􆿳��q'�vqng��#:�LH�ҋX�����jƓ�[���Eu ]����b3�'���Xw���\���]~'�H��{l�f|��rs�i��s�٭�`�̳��i;�������T�\ ��׃X�"��⹌y��o��C!T*Y�{'%s�Ǹ2���_�A.��vV�v��g��U-�eVJ:�~�ĬS�V���<��z��}�\w��0]~�ӵ(r7����b3�'���Xw�j�7������}0`a(􆿳��3pCtA 8�����;��]�JڒLy�]q�I���;E�@���=�tK �_"p��W�W��<��W{0`��!�6qK �_"p�{nr���<��W{0`��!�6q��T�Ѓ�Fu�%r�=y�"w߻Yg�����w�-�L��m+)q����h��@:S,���<C���O�G�}�(C#ƀ��=���a��bǬ�=�M^���B!.��@h�^fC��T�z���,}l#�mJ�0�6��������x�&��'�q�BZS[]N���B
��������So-�>�6C�(�HB�O�=��ܒ��Ek��[8{�n�_ �����p��Ss&	�&�
!�`�(i3�ݚ�Н���2�ͥ�lz\�Q��v�r��Rϻt<� ).�x��~\A�أ�g��~�	�7��7�ܥ��2�/��:M/�ա�^�jj��,}	f��J�/`0�����������}�(C#ƀ��=���a��JLm|��(�a��Tk@�0t�bGD@�F��qW��Ґ�Yj:{b6��P'	����t�\7�ܥ��2��yD�0Np�^���17T1���pY�~ȸDz�b9����$�n�����['Ȑ2��;�Q9�	d[�̮�U� ���_j0��.@.k���n��@��P���"5���q�؅��FJ��/��<Ӭ��['Ȑa:�$�77�}�(C#ƀ��=���a��JLm|�V��_�$2���w�"]W��n #�[��0F�s�ݺᣄ�I^Ɍ�|��yf{��������K70y�=`HV7�ܥ��2�/��:M/�CՐ3��F<@�Bcj;�J^��J�Y�"6��O\7�ܥ��2�/��:M/�CՐ3��F<@�Bcj;�J^��J�Y����ߠTq7�ܥ��2�/��:M/�CՐ3��F<�+�����R�:�%��X�B�l�2�vD���?a@!~�X����Ѵ���Z�����q�����P5��٪�N~����=���a��z>�n�S<�6�Q=�b��(��� �5�v��je���Yt	�����\�����!�`�(i3"�,�>E��4];ˍH��\�Mb�mOVy6RTsȸ�"rRY�<�"��@?P�Zv�!�`�(i3!�`�(i3 ���3�ҺIÙ=�H���mL�0ޥ0D���>M�J<0L�J��2���!�`�(i3!�`�(i3l0��F��j �i7�sp>KW℀4٬i�ۑ 55kU��!�`�(i3!�`�(i3!�`�(i3JHn��z��r9�3k��u���f�:X�T�f���y��̨!�`�(i3�E����F���8�TPm=_g}b��7ݲ���!�`�(i3�*���<�Hr�»�>��-U�f��Q��z�n��!�=�4e=��-	i�/B�6��&�elZ�_Hsȸ�"rR�%��ZJTD�l���tL!�`�(i3!�`�(i3 ���3�ҺIÙ=�H�<���͹W�D:���_�A.��W>����!�`�(i3!�`�(i3l0��F��jT�����NM��%�p@�R+��r