`timescale 1ns / 1ps
/////////////////////////////////////////////////////////////////////////////////
// �ļ����ԣ�		ģ���ļ�
// �ļ����ܣ�		��λ�źŲ���
// ��˾: 			�Ϻ���־ͨ�ż������޹�˾
// ����ʦ: 	   		XLX
// ��������:        2010��6��22�� 
// ģ����:    		Reset_Gen 
// ��Ŀ��:   		GNSS_Simulator
// Ŀ������: 		EP2C70F672C8
// ���߰汾:  		QII7.0
// ����汾��		V1.0
// �����ע: 
/////////////////////////////////////////////////////////////////////////////////

module Reset_Gen(
	clock,
	reset
    );
//////////////////////////////////////////////////////////////////////////////////
//�������IO���Ŷ���//
//////////////////////////////////////////////////////////////////////////////////
input										clock;
output										reset;
/*********************************************************************************/
/************************************����ο�ʼ***********************************/
/*********************************************************************************/	

//////////////////////////////////////////////////////////////////////////////////
//������λ�ź�//
//////////////////////////////////////////////////////////////////////////////////
reg		[9:0]								cnt_for_reset;
reg											reset;
	always @(posedge clock)
begin
	if(cnt_for_reset==800)
		begin
			cnt_for_reset  <= cnt_for_reset;
			reset				<= 1'b0;
		end
	else
		begin
			cnt_for_reset	<= cnt_for_reset + 1;
			reset				<= 1'b1;
		end
end	
/*********************************************************************************/
/************************************����ν���***********************************/
/*********************************************************************************/
endmodule