��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G0��@h ���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��:%��Z���xN��g�.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I+ĂiW,���D�+y[ف���rn��mo����/~.)��3�(����C�X��2�k(����)O��Ξ4�"�\�� ���K�O�{����a�s�Lj���ƶNc\֣�I��B���t��|U|�/֚m� �+d��.8%D.��n�P��<2�q�U��k�8u[\E���@N1�w�0XL����[fe�Hs��9lSUQ�S��)���2Ee�Y�R2
�I.��	���
����k�������0�?�}4��ѕ�������U��=>bMab�	;4��G����a�����(�I�?g�f�k%URPx�ζmR{z�W ���������	x]�fX�eϝ(�Я�mڍ'T����X�w{������:�%�+T%2q򋙔�M-US-�8<�n�У�Ǝ!�ѠV�>!�/�7��u���nEA��l���D�{��/Ƽ���\�4�sP	�b\qB�y$h��ݔf5*`]�|$ɋ��c�~�MUs c�+պNE��#Y��#p��'��������S�����:�֣I���Y/��S"�:����:�wl B����/��;��|B�6L����k�y.�)$����\�4�s���rH
>TT	q��$�2�����b��ǾI}`�~�MUs �?oQ�%'�s����o���_�xm7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3ts�JFAa��Bzb;ym��+a��ʁކ�+��T��C�NJ���1�:�Ω�*���g S)�-E�؟��%H�$��ī�o��<�)�G!�u�����!�M��E��c�W_QLuZoO�=���@$"��ea�8���*���g S)�-E��ri�y�!�3]o��in�m��+ r���7���?�_�K�E�\��Y�ea�;y� ����t����M��Ґ�m��[���b9����{oS�����\{F˯�+)��n̈́�zL͊�q���Vǃ����ܼ�Y�d5�:�wR�^Ƒ���b9�����%PM��NUkʽOy+W���F�^�g�&�0m�b9����s�AJL��؍��R��j�.(Wx*��|��pS���c,��-��%Mό���.��_F�k-�"�,�>E����-��%Mό���.ӳ�
�	?�<"�,�>E����-��%Mό���.�q�\E��0�����?x��#��]����������ݹ�0����9Cd���*�=��X��ʙ@E>*;�¬pX��g��U-�e�,���6+�\.�l���Yl���#�]�!��	Ǹ�y85�����5��d5�:�wR�^Ƒ����"X��[�'i�! ]���f�+��T�����h�6ؖ�(����C�-�nC/$������Ls�F�%ܪ���PL~΄gO�3f��*����"�Q:�{�1��q�©���ZO���]�(��0��r2���c�hm�i�]�׼�a�r��AR1<�N�؆�B��W+`�x�oP��@t�&�e�5
��Ib����rs�i�jf� l�Ǜ������CyW�f�tR�wX��}�
�?�?KYC'v���pG؍Y�]�׼�a�r��AR1<]Q�I����踫g(�r��3c���jj[}�@��Lr7�r��#[�f����0�]�8��jJ4P;�Q���n��̒��b�|��Ű�G�`��3�V2��J ���Bl)���;��q;
�Y5YqJH��[q�t��c_����+�˂߮<uw��˪?�-X��9cѶ��H�Ad�d��G&Tf���t�\~ �g8Yw�5�%]���a(􆿳��?ƾ��"}�`�W�Բ�������|����OxtX+�Y�z~~�Y_"R�W�u��"�A+�W��^�����f��|�F7�_���ɑ[�!�`�(i3e.��i�X�_�0��'nU�s��d�\;Tti��o���(��i7N�_�z*K�D�@�Y�4��j�O$� �;��|B/B�Â���P8��PS~��/��C[�[�l��a[�S��Y��Pv��?�(3z��z~~�Y_" �g8Yw���P�7� aT��3G?�d���&�*:W�q�qR7׷�:��ķc����,�p1ɠ�z�a�$��;q������it	�T���-M+��;��|BwI�u	�ogRr���R'cf���6�����m�F�!�_H^R�P:ض!!;��|B'O�d��FiI9�o�?�d���&��9�|���lm�����ȫ��=����t�����+�9�f�j�(� ���ָ�m�F�!�_H^R |~�($U*?�d���&��ݚ�Н�	9�rѮh�φ��<�6�@a� ���N����ݚ�Н����+�^U�	Y���;�jmT�#bs��2[�a��o���H�RtV�^Zt%��m&</)+?���Tif���GK7͍��|��W&":�ݚ�Н��̢k���"��w6�0��ɗ��zi#Y)M���Fe���2+m�7m�T��Ʈ+ˀa��z��2�,!�`�(i3e<�Ia��la��o���H�RtV�^!�`�(i3L�^��*�d�:��5c��M-03��N�L���Tw�f�H�;�7��w�@z�צ1�m+�D8!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �W?�;��M�S�"����}�ߗ�oHN��R��?�d���&�<�V�QK�}��C�Y�\�<�V�QK�}7���V�<� ��N�)gH}�BrJ�o�7��_�*
Ae���j���s��d���!i��'T���+�su�;�W6�o8:4�I���c�90�Ǘa��x�0�9&،�`����k��M�\���F�`yx�>�+X�M?��y�!�`�(i3FkH��۰H�J�������صW�my$�N��o�/���;!�`�(i3��$���͜P_�_S:g�RMm�o��'����Tj��^�G�E�BS�+��U�,�P!6���r����;�jmT�#�,l����M?��y�!�`�(i3Zt%��m&</)+?���Tif���GL�^��*�d8�˚��9�@�VҒm�!�`�(i3�5ߧE4��!�`�(i3��Ě�����}Dq�f��Fr��j&���"�g7�^�+:�I��)���W�w��fDIp��u���E�i�m}66j�"Hs,�A'��/>t.�66j�"Hs�@�6�_��V���(%����Z鎬�������(���q����"���0/ܤ�(g��V������Jƨ�Jt̫j(&
M�K;��%YM�	�v�3��3c���jj��8y�Ɋ����Z���F%�X�ԼQ�}�p�?��X9��ct�:��REs�N
�u�}�T�\ ��;��|B���r�����<��>�چ��n��r�v{��lw	�����?QZ���>$r�t�}iV��	��y�� �P�qN'Ds����V��	��y�2B��$�ij�}��VU�簦!N�'�y�G