��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G0��@h ���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�.�&ʺr����$l2�W�K��N<��;���Z��4d��{�
��|��Ȋ)zo1���á-�w~��dF��8�ĭ��Sɿ�{^��1�:�Ω�.�&ʺr����$l2�W�K��N<��;��� B]�pE���	x]̃Dj#^Da����M���v��W�&��v�=�z����)�,�˛D��w���旴4�����<��a��rl�ʩ{�Bf��QՊ(�
�d?t���raУ�Ν��u����l�|���j8��6�ܬl!����Y�f��a�Z��V���҂�L�?c�ĭ�t�k���er����$lkDP�%[B�o�O��XI���Wc"�b#Ӡe��?�F��&hWw�d�pP~��)%�����D��2E �c�=0N���6��H4�
� �AH�}��� �Ȱ��-+�T�8�hF�_!�>>��S�O1����h��]3�;���[=�%�
�R�+�hV�;/=�n;i���2_�q�JX�����@�>��+R���RL�a)=�y�~ ���������ߤ����Q�=�>�v�ֹY���8＀�L��q�Jp� ��g������a6���r<����}�a
��{0��d#��翑��HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A����2�P`��������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW�{b�2"���Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ��4Z��ʬ�ħƿ�9c�I�?g�f�Jm*)�m��+���qH�Ո4Z��ʬ�ئS��.V&��B֥�(����5��}�:���JŬ+��/�����,��B	hI�ˋ������Kp&�@���k�� ���3�ҺIÙ=�Hr��~-���I�R���F��c��Z��}��	�d�bzP#�-������4Q��#��w21�X��|�C#/<���q��!�u�ǭ��k��?��}��7Q�� +@����������'�=�OT���0�4z�S4ٗG�D:�]��H/!�S�av>�)'l:}��Q�Ȩ�+)	Y���
Ta�~�4�k�|L����ҭٕ!! �ָ3�o�:��o�Y�#�Ez��R�>}1�l+Tf]�i�#�l�-Px���H��U��p騥%�W,��{���7K��;������(�\���W/�������m��Z�
b�tU��֜��3��TG���PIÙ=�H0/�+Ύ��M���R��ӟ-��[7�d|���XP�����<��no#��٠R�^Ƒ���b9�����w9�ѷ��[MD|����a��'�-��띂ii�4];ˍH�P�(e�X�T}u��Q��L(\Ӧ�$�̎�)NC���)ҵ���]���>����C��ǩGY��-��%Mό���.ӳ�
�	?�<v�ј�"��Z鎬�������Ӊ*��y�7/����p���Z鎬����(��eظ���N:��e.��xu	���S8�/ #O�)R�^Ƒ����"X��[��Q[R�7�� ߌ�˕�(�
t��Y�{'%s���'����no#��٠R�^Ƒ����"X��[�'i�! ]���f�+��T����)�G�o���sp%r�M$�*�#�2��%�&���#�{�0;�}����\Ҧ�^���!�U��}�o���#�0��r2��dNI�,% e͉�Xkc�G���A�ڛr�z���*u�)�ʫ&*7=�3�J	��X�/ ��-�p=��Gm�o�j��`KL[�{W�g���F�i;�:U�v�3b��{"���,���"��y�xI�2^)b��@ŋ��5k.'C���Y�V������p�0ty�P���Պ�`^��3�J��\�v�w�?�b�>޼�\�vř9���=��\���.@A�-�]s�(_�<�� ��b�FP&����҅JHn��z���������x�&�F�]:��='����R��e%�2�ͼ���y�]�F�D�+�:�G�9�E᭗��_��&Yd&�j}!��n�͑��LK.I�:���3k��g1�e%�2����莇����_����~���i�x�k������y�"�V��q&=�a�7{�rN�cZ��t�������:(�����c8?-+eN�T�!f�GI(M���s�v��syu�s����g�r���3�a{��67�O0{����V������E�B?�$o��3k��g1���?Zkܼ����Ҳ�(����E�ߥq�X��WG ��EV�XK㈛�prj�r���3���*���!��
�j��TG�!;��WE�|���p8�<l%��Jh��AmY�f�aV6�$pap\7q߽n�������a�"��Y����:���2c����h�7�_��͑��LK.I�:���3k��g1�?�,t�J`�p�m����c8?-+eN�T�!f�GI(M���s����m�㛂���a�"�B���	��Id�����m��Fi#�ǩRq�Lu*���c8?-+eN#P�j2E�?��;*��ICm�5S ����'���o|k�Lbc¦�.��旵���!&[�x�R�"A��kT�׏�����Mj���;��D�2�7�?��i,��&lG�i��m�P�óM�˄No�M���MJJ�Y6�B�����6��-�=q�:�x�@u���h���D��uqIUe�JHn��z�c�����<�W�C%�����+.�ؙ�b�?ׄ/�LE �����\�v�n��l������}�v���Lj��f=�2f�o��"��U�[в��*�p6�!"d&���"\���.@A�-�]s�(_�<�� ��b�FP&����҅JHn��z�L�����"��cWN�Ψg��U-�eJҪ��D �bYu�c6L���@������LI�.��tA���ՔأͽgF"?Z�M����o���wu6�~sEz���O�� ݖF�Ut�\���t��ױE$��"�t�
��s��U;4l$'�_��F�5����A��T%��s�`��ޙe�勶1W�V�bSTG�!;��WE�|���rw�&�z<a��N� ��靤�}O�y�9�3����6���@�2���]]:�,�^�;��%YMYo.���1��Y[���U��%:����Vw�\�x`��:�c¦�.�������.�C�G�nD�t]<�LX��WG ��Z����e3�*���z���;�Aĳ�ޙe����;*��I�m�/
?A��kT��ࡔ 4�Ux��.��p3��Q�;uojr쇤��$w�ǌ�u�ݶdɑ�h��,�������L�@��e%�pV�>]ʄqL$CF[�S�٬�>�E��n
V~$9l�)(�BV�m^�?&�l�{�k�)��;*��I�m�/
?A��kT��ࡔ 4�Ux��.��p�G�B��uojr쇤��$w�ǌ4�04�jf�L��e�q�Lu*���c8?-+eN��#�"���|1Cv��E��
�9�����-���ʭ\r��$��"�t�
�W��]���y�"�V��q&=�a�7�����gP��U��%:O��E.�"-n��j�S����3k��g1��&.��8ݽE�c�t�W.�c�&��h�X~��6�='����R����\���o����z�F���Dܪ?EB�>�oj:�����GEV�X�d^�ϓ��23�Vw��šB)�Z����~D=�G�j�AmY�f�Ƙ�r��5ߧE4���]��	W���/�zU�=�����?H�
����Ѓ�I 1��6aa o�:�����)�x��.��p�Q�3'ζ#��"Z1�Sc�j H��2$%-���t��B�F�w��$�D-�;S5b	�?O��9�WE�|������'��ϩ��z4�g�Sc�j H��2$%-��u:Q��v�E��kUȔ�Ƃ�=89�8�^iPŲ�@���rah��cWN�Πd �^�z'Z�S�&�+E����A?L�����5 �x&A���0"�ͷj�Η@��Q���Pu��6~)ՄR*��uJ�7nd�����U���X��K�kH
�/�?����U<-���[J�ذ2����������W)Sc޺ #dִ��팒_�>c����� !(`���7��0<��>!�*� �`��U��_fI��'�{�"��}g�����zL͊�q��io2�&H��ݫ�Q�����6����r��1�Z���=�0x� Ĺ6NÌ	W�آ��A����bǆh���;�KAmY�f�
������'��E��T�
�rW��]��C Ln��S�W<����GRG��@ጀ�]�W�m��8���/�n��l����eew�˭�ߜ��}�+�0+�]4��ݪ��Ca��v.kr��(̥C5���?ׄ/�LQ�D��Ln��S�W�.�p�2�zgf�z�;qǙ�d��hw�к�&�@,F˯�+)�0x� Ĺ68y�%�v�T��7bE�g�;�b� �4�r6���K�TR"KJHn��z�L�����"���p+��+s�$�`��Z�n��[���Åޟ6eF���:&z�!A�������Ca��v.kr��(�k*���3��Q��)�N���%Ɩe�;����J>п�p=	�˳͠m�xW�J�H�[��'n�^0o�<:�W�_ĵn(���˧�0z�cUL�ݵj�<o�5�%]���a(􆿳��1�Q�/L��Hf�=jd�m=�L|Dt��	ZĞ�W+`�x�oP��@t�&�e�5
��������3I^�v�[�9q�Y�{'%s�rOw����A�T�g�v���>�֔ض1�Q�/L��W�Ͱ7阒|�6c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85�-�)�{�Z��s��R�wX�՜M�q�Z����Z�r�Y�}-�п� W��$0���>���˿������N���%Ɩh�����<���,Y#A�_�=�����w�_�2��K�TR"K�g��U-�e5��e6²��E��]�؀ǏU�e��FR���'S/�_wπ>@ �R��P�9J\�e
`�q���ʭ�O7}�»����Ck�MN�3�Q�D��̣����F�z�C���qg2�K?\?��~]l�*`Dg�8�Hk��|��-Wl���[w�4��<բ�]Z�Cď��/V�h}�L00:�g��U-�e(��w��x��-��U���T�\ ���|.�TӏR}���tE�U>�f&��'!msR��������ƃTrb�Jhf�|�Y$�h�ya�����aU�`�K-����16X{�"��}�u4��d�bR�wX����K�Q��2�b=��*Wؕf�*F���%��R��V愽��h}�L00:�g��U-�e5��e6²�T:���V�s��ҟ�s�(�X)󿥠&���Z02{�"��}�u4��d�bR�wX����K�Q��,����*Wؕf�*F���%��R��V愽��h}�L00:�g��U-�e5��e6²�T:���V�JG!2�|(�X)󿥠&���Z02{�"��}�u4��d�bR�wX����K�Qʘۥ<3� ����|e�7s�9���o��S8��A��H�cBh}�L00:�g��U-�e5��e6²[9Md��]�E0�+��зq8�Ј'���Xw�j�7��{�"��}ϻ�_���8���/�a'�<� \��2{U	fWgjZ������Q]� _�rs�i�ק)"�僁�cSS�b�YG���R�wX��1H��˧ݥ�BR"4c��h�W.�ۊY�7#�xI�/�6	�п�I7��-5��|�Of�K_��1B�&�P /r����$lR��A��Eg��g���O�O����E�V赊��r��'�Oy���6ʕ�Q��������/�m�S��j^mE[��Xv,T�� �Ac�N�A`~G��?.�#g�k���.���d��+���ÃI���c�90��q�	_����+�^�N���5��x�>�+X�M?��yЎ*vzwιx� �Q7���$=Q7l��C �Q��Y��-=���]	"e��0�U+�qbp@��m-�*��BҶ���X �Ac�N�An��톕�����z���nF���<�W�.�P��d�<*ok+Q�h'�Ȝx�5W ��̫(8��ɮe<�Ia��la��o���I���h�w��y�7/��i8i�+o{�"��}�u4��d�b�dh_��tC=�qإ����+L�����g�s��l�cu�a(􆿳�e�&���6qW�<���c����k��C �r������[�4�f,�8�|P�nkCf�$e��~h}�L00:C?�Q䨈y߉�m�$/X*F��c�D&����\��H��$�)�vx�"m_OP�@[�_zβrE��g�Hb��ȕR_�ڱA�e!�.�9�s��20��غ�7��y�7/��i8i�+ot�M��y���_L�H�lʇ��V@�?���'�@-�?$"�=��a����#ӗ�bJ�*ku���3l>��5<'�D���`�{o��T�-=���|Y[�q�ô@*�\�H�[��s����S�$~��HZ�UF��{κ��s�;��\(�3z�g��+˘\5�q�l;1Յ��iÍ�ф�A�xR ���J�QԢ��!�'��أͽgF"?���p+���"M�RZ�y��K�ݽ��������D5�|أͽgF"?���p+���"M�RZ�xkx U�_@���U���&0�]̽Cl�;��|B���8U�֝_�j�0=N;]%z���5��Z"��a�d�yH��}�Xv�9$[{^\�4h�fa(􆿳��D!G�$��ּ�9��@�m�۶-�Ez�?���e���l��c8?-+eN��`�6#'�c��=�t*V�M��nDŻ�&ǥ��?�d���&�fTpgZ���jp�6G�k.9Z����t�h��E�&�y+q
$�үe������hM��1o�l�P��~R��b�1��C���5�%]���a(􆿳��s��u�:㐀,R�*`Dg�8�Hk��|��x�6���k�5���5�m��'A>��"X��[�`�L�iցc�����M�~�B$X���V��	��y�W݅�#�f�b E���6j�"Hs^x6EoufQKg
�3�]φ��<�6�V�ҁGG�.Mm-;���c�Ì=f��Z�Qw�c4~Nr_�mS8<�n8.����b#"���l� ��V�I�Yo.���Pg�,ǐ��6�I�h�S-^^B;�֙�K�J���bd�T*Q�D���AƖX�y��pAS��4V}-�п� W��$0���>�����nR�N�o��nF���<�W�.�P��c3�fF�5.]���m+�cq
��T���xvW'��}�3���cD0�ʂ�j�Ï��	�l�lM�3 �[�{3^��=�O�-v�*_�mS8<�n�܅+���2W������|��RCc��P�)���i���\E�'����f	������"O��~��� <���,Y#Ao���wu6��pAS��4V}-�п� W��$0���>�����nR�N�o�y�<�J��}-�п� W��$0���>����15o�5�3���XE�ƃ�6�<Z)��obtBK�u�(�V�ܼ�.P�s�6m�����TS4�04�jf���F��O�<�P�����os�鮊��Q�d�
T�>�4:��φ��<�6����#�8��dȫw��[`0�x5��c�!{p85U��O�w��;D!�N}�m��{�,3�Hs8���l�E�a�x��c8?-+eN��`�6#�`�L�iֱg#�����[�Y�x1�ӉFAԢ�a\�����*��|>����n������� N��r*@��Mk�Hx�C#�K�"a��ُ�S�g�УJ/8��d�\(r����Ymd����Ԏ��.j�B�˝�,`Cd�p���z8�3q_҂T�q�G{����c�cSS�b�ԯ�J'>c�<c�9�Fs��u��Ifvi��a-6�Day�s������0��X{J\��$��ɤ&�U��f���L�ΪA��8�|P�nk�~����,M?��y��o<Z�L5s�"��=l&�c%=�)�a�x���2�b=��������W�6?���Ө��'�hiC���i���/A��4�z�X
3kZ�KQM���F$ޗk �4�r6�h}�L00:� ^M'���Cҷ��e��Z9��]���#�0�bM ?Z����rW��]��C ����X8��8���/����$����I�Y��G�j�>���/���k���cSS�b�E�0#�4j�T�\ ��k3�od><}����4�xȀ��D�[b%Ɨ�U�QU�k��Jd!IGc�{I��L�1p/-����n��I�8���$����I�Y��G�����zyN'�a[μ3z� �z�E��M'�b�	�)�.�ij0���!{�"��}n�m!t%qa(􆿳��ύ�>� ']v1�_ُ�_��^��{��|M1�9$[{^��o|����"X��[l-���}���W�6?���Ө��'�h/Q����ߝ��v�Y/�ܜ�������#oM.������\�vŅ��J���rw�&�z<a��r�����˓#���U�QU�k��Jd!IGc�{I��L�1p/-����n��I�8z�X
3kZ��<GHj-�_�r�� �W�6?��c�!{p85ˏ���|urw�&�z<a��r���+�uB;y��!/_�L�Z鎬�������(����#T��Ȓ��lXa-/`�z'��Ba����������w��o	�x$��@���E������pP��K:+>����YL���dȂ�Ͷ��.�X��WG ��hw�U�1�he�C�Hc�|��g;�X��WG ��d���T��jsrCm�kp�z����]v1�_ُ�_��^��56�6�ȃ'�)�Բc��bGW�A*k3�od><}����4h�Qf� �X��E=r5J�Ӝ$����b�Bϱ���2�b=�������AԢ�a\�	PcM�9S����q��k��\�v�07������"L?����o<Z�L5s�"��=l&�c%=�)�a�x���2�b=��������W�6?���Ө��'�hiC���i����  w��_z�X
3kZ�KQM�����$��P"G�wk�]���#�0����x �a���=7�I�Y��G�����zyN'�a[μ3z� �z�Ec�}���Fo|k�LbB�R���>_d���T��jsrCm�kp�z����]v1�_ُ�_��^������_M�<TC�}�����:(���27:����aٔ^?�����zyN���:��KY׏�����M'Ƶ�s]0{ɽ��&k@C�Ɨ0z�cUL��.�^�,��K�$�z�X
3kZ�ڱA�e!�.��t�>/�u��,P���_Wōd>A�T�g�v��o
���^��5ߧE4��
��T���x�;	㯰�$�)�vx)�K���'�#�c����ҷ�R�Ճ������-��U���u霴ԭg���NBq�`c�!1 ��Ktf*�gLYR!�rE�j��8�b���=+��<��](�!���`���\{ف(�7���n��T����C ����P����=�WK=Z�R�ڠa�r�"�R㬽�mV2i��h}�L00:�^Y�`��O7}�»Z}�R+�!�'��أͽgF"?LO��M|�sPn&��|�"���>� ����G�e� U_9^���\�}����� ��$A"u��p$(���%����H���=磡��{��1Y�[�2(���($�|�*��=| �����a��Y� ��|����:�����A�A�C��-eh�/�Lg�c�!{p85/Q����ߝ��vԩ �E�p�g��U-�e"�A��"�Y�{'%s�.W�jb��w�I����؀ǏU�e��FR���'S/�_wπ>)}���dG3;�hs���p+������)O�g��U-�e���+s�K������W\�y-T�OB �4�r6�h}�L00:Rl�I~�/T�K�^d��]�!��	Ǹ�y85���H�=fG/�'8k�{��|M1�9$[{^��o|����"X��[˹�H٫!ԵưT҃�1B�'�7�=;v8�^�W�U����*���/Td@��c�����M�~�%�,�х��J���'��������_(��R�#�"-��K�TR"K��L ����r\ڄ7
�?�d���&�use�	��EzQ8�_53r�Ny�v��i]�>�u5�D��7d��c����P"G�wk�M/w����?z�Kv��oV<��/���^�:gʶ�7��i0�n��ϵ!�f�G�y-T�OB �4�r6��cU�tFZQDu����-�Vb� �Z鎬�������(�����I :㐀,R�*`Dg�8�Hk��|��!�x�����!�=�ߝ��vԩ �E�p��"X��[˹�H٫!�M�0���j�>���/���k���cSS�b�p�[k����Cҷ��e̷_��yC��S8�k��m�ݧ�G�y����k�)�;�,�m�۶<��%��������O%WJB8�^C
�6n�$ٿr�Ի;_W��(ξv�釰G/�'8k���3�c����E����P�++�hW�w��fDkL�@��9�GKP���hG�*	�B&hL��C������Q5r�����#>�;��kh}�L00:u���Y`i�c�N��j��n<�s��;#6ʮ��Vy���Z@�05޳�˚��i��I���PJ���9�43Iz6k�c��2�b=�]��E/y4����ןw<LC9s�� ���c��Ok����R�#�"-h}�L00:;��|BqR�ϵ�i��,F�d�h\.;��L�O���X;����C ��kT�q�!D�t
��5Zbz�Z�f�x�HZ��,e"75�EZ��s��rN��t"O]��!���c�A�L'@fU�X?0I"�`�it�M��f�֝_�j�0=N;]%z���5��Z"�'��G�<���,Y#A	u�e�2�?�m�۶�so����O7}�»�QNȮ���k/��m#�J'�!���=�@q��u���"6ޭ<:�&.am� W�����H��6�Br���N%'tF��;���R��C� �Y��#_1�|.�~� �����$�\՛��2�k�S�{ �d�*��M�,4#�rQ��G�t>��Kò����{��|M1�9$[{^��o|�Ψg��U-�e"�A��"�Y�{'%s�.W�jb�ԡ*
T��Õ���PLJ�/���k���cSS�b�E�0#�4j�T�\ ���O�����7F1�	�A
�)�𭅐t��PЕ���PLJ�/���k���cSS�b��6N|���ʸ��g?��f+��hg�grYn�9�f�u��L;Ӂc�����M�~�Y�5� a��2�����Vc�{b�'���Lx�ƺ�M���	�n��XU���#fhr��y�ڔ�.������������/�LBgh�c,q������z�.���f%%eo���sp%�j����P"G�wk��%R[�]db6ڏ� �7.�O��S}o�"_�cSS�b垊*��䮻E�&�y+��2�b=��E���s��U��֜��3�T�\ �͊�51�X�c�rs�i��]S���D[�l��a[�S���}o]�
\j}�C���&��vt�*��]�3���p+���b"u2��O�/���k��Q�D�䀭�ĭ��Xw��l(�i�g��U-�e@�0Iݥ�Mj�(ȅ��Z������ܓ���'Ս��"���<'X�|��I~�v�(�>�{��D�h\�J���/�hD({ՒD�jט~���@�5�^R�[ZD���Sd�o�#���Ik�m�Q�<��W�2�ý������W\�y-T�OB �4�r6�h}�L00:� ^M'���Cҷ��e9f2Pih{`r���	� �4�r6�h}�L00:� ^M'���`y����p��*
{+Y���>�[6: �|J��q�}��k�)�;�,�m�۶<��%����'�]C~�̄��v���&�?���B�+�V�p�nB�W��`6j�"Hs�MSYQ
�m1�H���W�w��fD���oaDU�KF��J���64� �Ac�N�A Ҳ́p��xkx U�_@j`���؟�1�:�Ω�����|"�W~���vْl��]�B�7's0ۉO�?�^"��@���k��!�`�(i3����Oo|	J�^�l��?��X{yAuޞ�����i���a�����Օ��qvdЧ^{�j ���X!�4V�H�%p"��RfC` ��\U9����u��B�bq��2*Q=F�k�mD#V��[��"|�W������Ϧ^c!�6 �ef�/EI���ā4@Q�/�`u_=3O�̃苇��Fe�.��=")r���ꀍ�˺�Q�����+�+:��M���ʦ�<��K_�0ß\iygҟ�%ў׫�Jd!IG�,e"75�E��W��_�ړ8���/��vsi�����zgm##��+?B�OA4�G�1�/�;�¬pX��g��U-�e�kH����V��	��y��dm����a�m��W�^�B�a#���l���Z\��C ����P������)T�FdT���+��@-�-'͏����������ܩ�x�l��1�U� �1�}�W7��c�r��]n��-��M��lU �Ac�N�A��8&�N̕�;}��)�[���6�X;p`�h�5,Wlr�r%)cAI�x�~����4��)+�[Z��?d��A �4<��!I��X��$�� 9Km!Қ��B����3�=����m��:r��gx�n�W�����v�o^{�����O,8�֐�f�-�X;p`�lsσw�kzU`��W�.t�%�Z?��m�CY���:��ZEG*w��qĝ�&�����B�_����4,�Q��{��|M1�9$[{^��o|����"X��[֗Q"t����x�Jma,���^��5����PLJ�/���k���cSS�b�E�0#�4j�T�\ �ͮ$CqaEW;6j�"Hsϣ%�?��s�z%�ژ�(�2��Ȅ&N+e���ٿLv�$�`K�'$vr�����&�j�^*zV�}zj>gm�$�kT
���ۚʦ�9b	J?QW����h}�L00:;��|B�����Ղ}C&�Cz�m�۶<��%����=<R��ޟ�����'��Y3���6�AmY�f���=����E�VmM��}-�п� W��$0���>����_��nk�kB�:'���e2�%V��J!��m�۶<��%��������O%WR�wX�չ�G�Ȧj�E��g�Hb���FtY�����|�wc�e9��%�+ Ixcw���Z�����~���I�����_�9$[{^��o|�ΰE5CN%�Z%����S�v�b�kA�T�g�v��^��r��1�R��j}�C���&��vt�*��]�3{�"��}�}P�.{��|M1�9$[{^��o|����"X��[�`�L�i֜���,�ǰL�[��V���Z���V��	��y�f���{1��c�ҩƮ�Jj�'de]�3{<�Yo.����-��U��?�d���&�Tx(C�����D5�|أͽgF"?{�"��}E�:]���A^���\�}�DѥGu��0�]̽Cl�;��|B��mi׮�N�[��|������hM��1o�l�P��~R��b�	u�e�2�?�m�۶<��%�����"�S��rN��t"O]���q�}��X���4)��m�۶<��%�����"�S��R�wX���P�++�hW�w��fDK�R����d�Sse5�U>�f&��'!msR������O�[(`q�}w"�5 �Ac�N�A�a�sL�g��U-�e;d9ךp8�^�W�U�}w"�5 �Ac�N�A�a�sL�g��U-�e�SB�9�H��L�%��x�-
�΁#g�k����ξ�|��U>�f&��'!msR�����נp�Qe�L�����*����6��	���Cҷ��e�|��*��U>�f&��'!msR�����׽��9\�	Z���/:���lC��U�T�\ �ͭNjX�U�6j�"Hs�x�ʤ�^m1�H���W�w��fDP������@[�_zβrQ�ͼ����b�A`�Ҭ����5A���t�T��S�,9!:-I/B޾Pk���e��q�w~��A(�c���_G��Hb�ñ ��3�JJݾ�'�\{ف(�7��<�h�#���C �AƖX�y���?~f|��d�����w�⽒�;��c���XL;jy"k�{H�3)-)��m���� iJa��������ܖA���ol��t;N�09h\dN�<@Iv��nt=:ྵp�!����&^��b5�sw��
�(�V�ܼ�.�%Υb3S6 -�&���^a�nu4Bޗ��jw�	��-��@�%rk�,l����M?��y�NM���������[V��M*;��c���X�8vw��^C\E�'����f	������"O����n��T����C ���Ǭ����RO�?��~]l�*`Dg�8�Hk��|��!�x�����_|���N�[��|������hM��1o�l�P��~R��b��N*�95��{b��vW'��}�D�Tu�^?�&^��9�׍�����u���?�)����^�{"}W;��ܐ�}�۪�G���_��e0�@\}p