��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G0��@h ���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��k�	G���%��%���UQ���?6U���T��ײ2��>���^k�/7�?1�(�c��ly[�$D֍r�	�tX�)�`���$��[dm��+@ˏ^ow�Vx���_>{������6��H4ٳ�k.w�.u���ŏ|{T%�at�3������ͧpJw �^���Us�JG�DGsc2�aB�>�;�C�l���o �����$[Z�i��%A�a��gs|�e
�9��Ax!P����9SA����q�HS�b"L]$7!����Y�f��a�Z��V2 �Q[7U�i�#!����P�>ol[�y������{S�O��<$e|����w'��1�:�Ω��k�	G���%��%���UQ���?6U���T�����\�4�sP	�b\qB�y$h��2���[emدQ�s�u�5Q�o�FS��n� F{�B*�2����_]�
K��&Tj�P�6
� �AH� K�`A���vJ�^��K+¬�I	�_�Մ�ѕ�������%"�;���
r[��<h$p<��|�	���k�8���҆�|n���:�o�E��ĕ��(�$��W��ih ��ѕ���Ϫ+2���O'{���O0�UxX�1��J'H��q�k��Y�"�+`VU���`�+N/��Fh�a~��1���VY�x��;K�:n##���Ψ�	�ǳ����c,>0�~G�6�&�^C��������{�;¬>P�2-i_��2f¬Y��RL�a)�O��u����H7�'*�O��3Q=b���{!�zg�Z�$gZߌ��h}�0�iH��L�8$�+:H뉉�V��=ƨ7K8� c��(�U����	x]̍��;��+e>�� 6V���~w���I
>��������V���8e3Z}�ax�� 5���_�xm7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3ts�JFAa��Bzb;ym��+a��ʁކ�+��T��C�NJ���1�:�Ω�*���g S)�-E��ri�y�!�3]o��in�m��+�<4��ˌ�ň��h���T�%�/ң��n�
8JAZ�NCIw4t�iZ]XF�������̇��� +��u*K6HT�����Np�S�q����E©�ʐx�?�'n�^0ov	��ě�e>����C8�����M�g����"�,�>E����-��%Mό���.���|��pe���b���|g�Y�'���Xw-�}��dӅ� T���c��Et�Y�{'%s�:�f~=g(���B���o��+eQ�s����|#9���>��682�6�d�fc��Et��q���U�[��N�������l|���(Z鎬�����
��al>�dN�0F^�S�����5	���]���c�A�L' �oy�
!��9b�S� 7�v�ԯ��Q[R�7�%t̓�@�3��ra�ʄ�TD��ό���.Ӂ��̰�!)����bX��|g�Y�'���Xw��E�d����'(��Yl���#�]�!����M[��Ǣ=�?��3�*�p���@IE�U��>��l%i�-�%t̓�@����9�T�TD���rs�i�jf� l��E�4.@�7��y%%\�HP@�a�~�7���� ��JL�N{a�9Ow�Y��k��ı����V���}����W*�׸-�nC/$����[5`� Oag�qod�֓��+��T���jB�Fg�Y씤`��p}RQaI+اy�TՄL�Y�͋�<��P�x��r��VYW\�'g`$�Y1#��Z�����XP�����w�K��ݑ�][H���\Q^���0a=cj<���|0���)ÒPl질�z���	_=���CA9�9�|�U�m�l��'�5�e`��9nS�dB��,�:U�h���<��j����k��#�M/*�3���+��q2/��q�&��DP֞ �'��L�� ���3�Һ�cY�~�"���ʷ������<ҡ��~d�O����������P}�2�H�uv*@^7&ģMa(􆿳��ȡp��'���Xw�j�7����'�\�n`��!��B�T�\ ��Z��| �ƐkѶ���� �(�Mz�Iʬ�v�z��]��G~�Ϲ��T䘚�C�h\K�5~�Wv�A��2���HF3}�
�?��(R\֎u�eK�	�$V��d�٣���N N�S���c��:KYЙMǿI?��u�Op'���Xw��
IǬ�qcW�(u�" Oag�֠$b#^M�Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�ˊt��q���1U��3{@�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc6^-Yu�%�n��UM>8c<�@�׀%5F���>&S�XQ�� ��&�>&S�XQ���<�T���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�fYCJdR>IE�ث㭕�K��ShO��7�� ���ѡm>OM�Ѫ��z4�֏`N%�W��J�� �.4%,��ʇf�Y�����!>�j�V!*2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�C�9�*Q����t�T��?E-h��`f���sd�G}%����3fJX ����X��S�Ȓ�'ž1�|�'�����j��c�Q����̰�!�Xy|�W�#QSU:��8���[{/;k+Q�h'�Ȝx�5W ��̫(�H��
J��͒t�]��/",oMG~�>y�pA��x��w�����$J�L߉���v�_ej�x@3��0������0��G���_��b~*��s��(R\֎u��Gj7�uz�Va�ir��[��o}�N���Npu��r�偘�̰�!�Xy|�W���d�L����|e"��jVѭ@��l�^!ЙMǿI?v�h�C��/��kOT$f��_Ub��7��G_���;�P�t�5�׹�_S���\���Qw� q���`p�~(�M6����Z9��	h��4������l�Hv:g7���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�
t�������t�T��?E-h��$^(?��"]�B���[�.��|ȃ�A(�c���_G��Hb� h�ҩ�q�� �����e���߆�p�h��d��JXl'�T��~��Uг�|<�#�-�p�g2�I�7����_j���?\�z?Xk��;�P�t�5�׹��ܜr�a��t����=�Y��q�$���t�T�z�����#�ɼ�ϒ�����^����ܐ�����?)zni�յ[+8��^�鄃�ջ^B�}u��ݓ�W������E����3��Y$�VZ�ڋ���Y���u��T����l��M��/,;�.��1���-����!�`�(i3��w�`L�U5���M���[ӝ��o7fĉ>99��j���GpG�&ց�*�^rPk�`����>e�FW�DVx>74/������������l��M��/,;�.��1���-����!�`�(i3��;��L���W��7=G��Hb� h�ҩ�9��n�7�Y���_j����[�SRC����P�Jb՝� s�#���k$ 9��n�7�Y���_j����[�SRC.��:����%>�rGO�D mWN՝� s�#r%�:e�q���f�e�&�U��f�!�`�(i3oв%u�K����^���'ƃ�3�Y1tSjv�!�`�(i3����-J݉�|�T����
�:qEp�;�P�t�5
�:qEp�;�P�t�5���aR��ݓ�W���s�U����&U�)j�S���ܚ��@��f�\%����(�̚�ݚ�Н��"� ��.q���f�e�M?��y�!�`�(i3oв%u�K����^���'ƃ�3�Y1tSjv�!�`�(i3����-J2�բU�?j���4(!�`�(i31���~!�`�(i3����-J2�բU�?���~t�!�`�(i3�5ߧE4��!�`�(i3��Rx��íN=]8k��.ͥ�H�RtV�^��#�a�Ą��$J�L�l:�
d��>��(��Z!�`�(i3���ܚ��@��f�\%���M,�ݚ�Н��Ra])n#���r����!�`�(i3��w�`L�U5���M�����yV�a{
�:qEp�;�P�t�5
�:qEp�;�P�t�5���aR��ݓ�W����q��F��&U�)j�S���ܚ��@��f�\%��	�3���ݚ�Н��"� ��.q���f�e�M?��y�!�`�(i3�H�?��颢l��<_9}�	�-�ud�����b/?�-NER�ڵq`�8�I�Jh�Ġ�Ǟ��3��T�DF�W �!�`�(i3��Vb�#�9��|���׊EaP���n����7���yꐳ$�(�����k��
�~yj9�?�Ȏ��$73�!	�Ø�e�!�`�(i3��Rx��íN=]8k��.ͥ�H�RtV�^��#�a�Ą��$J�L�l:�
d��>��(��Z!�`�(i3���ܚ��@��f�\%����(�̚�ݚ�Н��Ra])n#���r����!�`�(i3��w�`L�U5���M��4O���a��
�:qEp�;�P�t�5
�:qEp�;�P�t�5���aR��ݓ�W���	�N�M��/�9ސtjCH�d*��=����h���>��[V�ݚ�Н�;�V&S�b�4���n��Fr��jL��[�)�jMO����i���q��:�Պ:�a���%t̓�@��5)��Z^�h��N�M��||�r !$��=m�n��z�w��"�on�tUk�.Ot��[��o}�nqY���1���~!�`�(i3!�`�(i3�>d�g�K���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ږj��Y��f(����#�f�45L���.PyBPȥ�BR�����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ڧ�wFB�b���t�T��?E-h��`f���sd�G}%����3f�F�f�V�2�~ڦ'ž1�|�'�����j��c�Q�;�~��-�f����Ga��'DV���b�z'hۉ)K7͍���E@���!��"� +}0�ʂ�j�Ï��	�l�lM�3 ԫ[=�.n�9�F ��T�#"c���]��&Y��V��|#HK���V�,��8�Eʨ�`N/�<<��lp��N�DNl�'}����=��,:&�fh��[�? ���Oρ!�`�(i3�*����;�.��1�](g���М��^���'ƃ�3�Y�}	Vӯ)������7�	��c��*!�`�(i3�r��f3K����H������P��l_��H�Ra])n#��;��L���W��7=#o�]�ʄǬ�$gQy�f�[����U1tSjv�����l��(�Mz�I�ݾ����]2�lـ۞���v������#{�$f��_Ub�F�S�1 �ї��Yt���:!���ԫ�o�u�/]ƄWYH��\!�U��0�|섃Va�iryP��C��?�T'�����|�x@�"�onq�.F'��_H�RtV�^;�~��-�f����Ga�\�׺h��I� �����ݚ�Н��5ߧE4��HN��R���ء�I��߸��S�Ȍٽt� $�N�;}it��j�3��ԩ v������b���%w�*�7��quA0�e]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7���_J��`��Q�����7�癆cgQw�c4~Nr_�mS8<�n)�{6�U���(R\֎u�J�
�M�K7͍��|��W&":����@|����^a�nu4Bޗ��jw�	���k��M����c!�}q���f�e�x��w����ϭO�cX.��m�T{
�z���=�9��|���#o�]�ʄ�;4�zu%��XW�G�<b~*��s�
�IӜ�_���ˋ1tSjv�ݑ���&�dh����Mԓ?��۳lU`7�X��=�̢k����(R\֎u��Gj7�uz�Va�ir�3i��U��[�ܡI'S��0~�$֚e:(L����-������l�^!�%��ږ���⣮`4hz�<Ρ��nh�"Mfĉ>99��A0ok�����F��O�\E�W��4b�^�#�nish�Ž���D��d���(R\֎u�ַ�����ڥ����Ⱦ�c�r%�乍���Tj'{w#/ B!�`�(i3?Q�@X>#��`p�~(�M�f%����M�{�|Lɗh�5��
�4���｝�b�Bϱ��LU=���`����ݚ�Н�!�`�(i3�>d�g�K{U��������pG`���IX0F�MV�ҁGG�.Mm-;�d=��¾ȼ\���F�`yx�>�+X�M?��y��2��}���'��L��K� |�>��̢k���F�KD�Vr[/}>5��0�B� �b���H��������0��G���_��b~*��s��(R\֎u��Gj7�uz_�mS8<�n�ݚ�Н��;�%�R���XƤ5_�P"G�wk��呞HXx�Ir��͕� h�ҩ�?V��j�c ��b;�^օ?D^��՝� s�#���k$ ?V��j�c ��b;� ,��rQob.�Y�2W>������$f��_Ub�F�S�1 ����F��O�}�	76�&�j���Gp��ܐ�}�	aF�oN��n={�ϒ�ք� =m/4@�s Oag�=ʰ�E�c