��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G0��@h ���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	��q5.A��|�H����VM.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I+ĂiW,���D�+y_�L_H��-..i=?�m��+�<4��ˌ��|��v��ӳ��$Fe@���N�w	*D���y&�f��+K��[y��ڂb�nP	�'~�c�:��/lt�3� P�;��1�-���f񻲗��~o��:���F�q�\�7Y[���G���d�֗r�5�c$e
�9��Ax!P�������H3����^�CG�1 T�V	�tL��	�<�A�}Q��	����<5�T7y;��S���4B�@T�,�찱�y�Zk���fi���60��g��b#Ӡe��?�F��&k�ZV"��s��;#�A�v�N<��;���u��w)�S�5� ��~篟|�<8�F�-:��ԧN��78�:r&@��$�9��_,n׎ ��73��>g�����Mp᫼���hvK+�va��2鍔�	g\A`�6��{���9��m�!=�y����h�}Y��݅ 0�����\���>k�"�o?�M��;]�=��)�I��)܅��J�|(�����	x]̍��;�������]e
X��r���Hߵg���jR�"�H�ٳ,�M(F�N��d�>�l;��r�O��C��0��$�>��w��z�!%���1Ѵl���u���;���	tR�\�Σ�cV�Y$�S�in���:��M�� B�h2�����{�;¬>P�2-i_ϐc\�sdHF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�����ga�^?u��v��[���y�URc���Y�{'%s��c2]�l���gZl�B�����|�$RqF���{��/)̡<�[
�=Pn��tw:g+��T��d^��_|��3g�ݜ��s8[Z�`
5��*�z�������D���J7"~����d��KJ(𬍝��;{g�P�r�|A�"C��dKBE�	g�yߓ����<�m��+��$|��;D���J7"~����d
��A�aG�+��T�����h�6ؖ�{��^�
r��4�3dY�-�nC/$jQ߰�H�M��RV!�`�(i3U��֜��3����C��n����e;��}Dq�f�S^�1���yد�9����)h����M��%�p@��\ NhJ���/�UI��?X�c"`.� �#�i0�[X�b\gA�[3�.!�`�(i3�=��?Q���n�;�X_y�F�!�`�(i3�{d��L����Oq0}�+�]}wӭ����?�+,���iVA�ڦ�c4���^���.�c��><�$�z�)
ԏ�.T٢ߡ[�1�g�=��2U�u�H
(����7S��Ro8�ih���
�e�~w�!�`�(i3!�`�(i3!�`�(i3!�`�(i35K�,<J��.� �#�i�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3ԁ�42����t|��z�W87"�o��ѾJJ�����	.l�@{���e����P];�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�-��\���7ȡ�/�!ҔkmB����I��%�)��!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=�����-VL(;�D��g�FBZbQH8�I�we3��r^�����!�`�(i3!�`�(i3!�`�(i3!�`�(i3m�z��P���ڞ��3*�f՗h�Vdoq�M辙�
so��j�!�`�(i3!�`�(i3!�`�(i3!�`�(i3MX����C���7}�jA�� <LS�ʌ���p5B���� �o�X�S��Ǵ��BE���Kt�I�ZMz��v�N`Z�NYUO��z�W87"�o�j'��y�?&�2�����B�X
d�E U�V|���hy�|�ր9�j���B���7�F����|��p+E��%>zcbp��'��}Dq�f�4��d�X��H���z{<���낌״$(�>g�!�`�(i3)�{6�U����/��w�=�J�5x������l����4�n���xǊ��T�3,R�^Ƒ�ӳt&:���aCPW�����8fDs;ly��\%�0�9&،{"�Lެ�k<�Lơ��*T�Z|{�0z�cULD�vO��|��!��5:A�8���/�l|�*"k���(ӈ���m�r�������Ȋ�?�Qs5��uYl���#Kv���:1�#���FT����fK6�L+�.8%�����dN�<@Iv��nt=:�rl��7�L�{	�����Wm�0b��"B��$%eqq�\L$�����//��kOTm�ڨ�hծ<�6�Q=a��	�sǡ �w�;>cbp��'@
9��yž
�I�>y�t&:���aCPW�����8fDs;ly��\%���y��lDJ�z`_�z^9;����l����4�e�kzP��}Dq�f�)�{6�U������ł�me":l�n(��̓iq�����f-���bX+D���0�7a
��r��X~L��U���N���{_8�Y��n3��v2!�`�(i3�ǽbI�͎DX��,�6�HaDl��+BY��9�)(����������qϛ�M~!�`�(i3�ˇ�h��]�Hlu�����}Dq�f�4ﲐ�if���ٷ����
t��{<���낌)P<�ܓ�Y��'T���+\��.��4��!%���Kv���ft�s� uƍ2���l�A�����2>�>���v�|��z'���Xw�����C��ݚ�Н����v�gY�����Iꑤߎ��J���T���b+}y[���S�fh�����0�T<9 =��9�j���B]��>��y�(�Tl��z^9/�~��e:[e��mea�8���s8�R�	��q5.A��|d,-��~7�f[l	E�^1pK���}|��QQ)������Yk"1/�<4��ˌ��|��v�����i9���(��j�:�`�@��i�+�.$X�j��Y+�K��Q�q�v�1��+N��2�g�-�:J~�n�E�T\�HP�<���^��k��K�+EC�����6��lC��U7�C��zC@Mw�Y	��D���F����dZ�'%�H���	8D? ʞ����H� }��D7ѡI4М_���ބ6cbp��'�6i����uٓ��������<���� )p�P���/�@����gGL�%�X�0g��D���p�VU��Jm�QA�Q* }�
�?�J-ڦ�.�5C�V���3��d�٣��c�A�L'W����I�7���&�_��lC��U�T�\ �͘�f��p�b�z'hۉ)��d�7�qĠ�B�D�F ��4 >y�;o�� ���d�٣��c�A�L'�����CyW�f�t��ł�!r�dN�<@Iv��nt=:�`��K Y�o�$C�J�ol�9pO�ڹ��1w�Z�>)���'vX[���U��m�Q G�f0�k�p�m~|��V4��������v.7a
��r��}8���uӜk��(���B���j'��y�?DNf���it4�/�7������k�tk���P����ڷe�cb!��u���p>�:�6Gި���Zu|]!T����ZBi�mR!.<ή�$*X�Ɋ� ����t���L	k���!qmX}���ZBi�mR�o��3�v����1؜��I�}jTc��փ�����k��zc�Э��8��d@y8��I�ע�s�B>>�W�#�y��7S��ZNV�n��`Ы��S�$�E�#s�8F`�K�;��:�~A��7Av3س��+K����Q�"x.2|Tb�f��zV�����[�#�؅z����T�K��`�/�.	Ѝ3!�`�(i3%��!�7q���Y� ���Ja���d����3&�.C������٫Np�a%��w�4	A�܊�k����h�Ӭ~[6���x1�~g_!�`�(i3!�`�(i3!�`�(i3!�`�(i3�c�n��X�n}?C�cU���?*����!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3":�=�/+T����c�~)�8![L~C�RpЖ�!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD�U �l�2�C�����������!����,=�p�,y4�N_��ʥ��ԩO�j���Gp��ܐ�}�г*O�v�mW��q?�� �U��C�^�D��&V��ң�O�?Q�8��I�ע�s�B>��vXٙZð��T�ݚ�Н�c�@�����.b�����2	�� �6�B��~5ʈy�@ҕɗ��zi#l�%�[��(-M�O��~�'E>�����Y��z��SͲp�����x(�i��/R<��}�u�4����&�)φ5e�+ż٧����D�d
 � v�)���6J��O�j}�8��:�x�05�2���H�RtV�^����K�}�7Ԝ7(u�/�"����1����߾��lP�#Ty�W1��X/��kOT�I���`��O�/=1>,Z3���ƍ2���l�`���*1�H�����ǽbI���.d�i�>1tSjv���'T���+�N_��ʥ� ���-�ݚ�Н���jVѭ@!�`�(i3��򴏓�	ܿ�B�MҜ�}Dq�f���Ě�����}Dq�f��ӷ�R��&U�)j�S���߂l��״$(�>g���'T���+��k� vpų���2zG�_h�����l���`�9<'�/�.d�i�>1tSjv���'T���+�N_��ʥ���Y� �>��������w�w:�!�`�(i3a+kb�Ϫ��Y��[�P@�m�T���%>�rG�@�	����ʁ���Mյ$��Q��@&U�)j�S
��X���W��Pw-��!~f�{���%>�rG�4���n��Fr��ja�U�ے
'E�=`�M
xM�v.����V�8�|��k���u&kA�-7�,���X�ޅ�S�J\7��1r��_dW�����V���%jL]�T!R͋ݗƩ���=�����@Ã�D譸nٶnڹ����|e"�#M�#/g�%��v���|#HK��JZ��=�)_�mS8<�n�ݚ�Н�z��SͲ����E�EqLt��.�Ra])n#���r�����B�G�.�W��Pw-w���nNH���%>�rGO�D mWN
L	�\k]�ܿ�87�ou����]_�m�tkK��?D�8��`E��+��'�^����J��N0�;�jmT�#�Ȑ�TA��M?��y�!�`�(i3�L	k���Y��[�P@�m�T�	��x��ݚ�Н�z��SͲ����E�EczUEg�>fĉ>99�񗺻�C��mJ�0�6�(*�O�qe��0�UMxw��f���W��Pw-��!~f�{HN��R��@"�����߸��S�Ȍ����P,���7�	寁��Q��o�mH��U�����k��zc�Э��8��d@y�Fq(�Kǰ�!f� �T$"��M?��y��
�*�ݡK�+���w����O״�b�z'hۉ)��d�7�q��H	EJF�d� �n�w��a�E�Rq���my$�N��o�/���;i�Q���d��i��7�����h�ura$�>�u�:�>��u��r��ϴM�ԕṅ ,�X6ae�Ɵ�s��H�RtV�^m����'K�j��=��\m����'K���uT�.�H	EJF�d� �n�w���;o�w$V%�kˣ����[9o�����5ߧE4����Ě������+Y��a�U�ے
�,�J�3�Ve��˅�ۊ�:�	�&v�5���4�ǽbI���}��u@:ft�� �yۂ�J1����-~J�
�M��ǽbI���}��u@:LKXkyP�%��.��^���L���1F�]�q:�q���8̷~y�Ys^�/+puhR�c�8m�ͣ����G���@&�>?DU`N'�[�	_6f�K0�FQ��ݢ��{� ���\�'%e��>��l�=��?qB2\�� �ǝ�,^aj�`�ud�kְ _;��i�1Yq�^Ȃ�	��LZ�K��V��?|����)м��$9h3bU�����%v�{�Q�^�V�)�:y^6gV���(��
�3[2�����Tqt���~��	��nٻsv�^��.��O�37�˱�5$�Ƣ�/몰���:qڅGÙ��܏C�;PU񩊭H�V������R���YƼ/E�g�������(ӈ��m���R��;��|B�0+x�@f��v!b�t5�U���~y�Ys^�M|�"D5�O�%E#P/8��A0�/ʍ�z�yL��n��p��b�Bϱ�m����'KN+?��T+D���0�7a
��r�"j���b7��I M^J7x��D���c�&ck����&FY��ښU:Q��V��	��y�s�|;�鞍��F ʔ��g ĳ
d�YB%��:ޜ9�6);��|B <�Az��'\��i��{_8�Y���˂lq��qgF���~�Ǵݵ��ح��tG<�, ����t��I[�=��?]9�(b���*5�����e����͠�)&�ܽK�+���w�D_Y�4�DUc�&ck���CyW�f�tR�wX�՜���,�ǰ��#x$E��r���c��J��N0�Pj�}|�^v-�b�+�