`timescale 1ns / 1ps
/////////////////////////////////////////////////////////////////////////////////
// �ļ����ԣ�		ģ���ļ�
// �ļ����ܣ�		AD����ģ��
// ��˾: 			�Ϻ���־ͨ�ż������޹�˾
// ����ʦ: 	   		XLX
// ��������:        2011��08��15�� 
// ģ����:    		DATA_LATCH 
// ��Ŀ��:   		MultiFunctionSampProc
// Ŀ������: 		EP2S60F1020I4
// ���߰汾:  		QII7.2
// ����汾��		V1.1
// �����ע: 
/////////////////////////////////////////////////////////////////////////////////
module	DATA_LATCH
(
	clk,
	datain,
	dataout
);
//////////////////////////////////////////////////////////////////////////////////
//�������IO���Ŷ���//
//////////////////////////////////////////////////////////////////////////////////
input											clk;
input		[11:0]								datain;
output reg	[11:0]								dataout;
/*********************************************************************************/
/************************************����ο�ʼ***********************************/
/*********************************************************************************/ 
	always @(negedge clk) 
begin
	dataout <= datain;
end
/*********************************************************************************/
/************************************����ν���***********************************/
/*********************************************************************************/                                                                                                                                                                                                                                                                                                                                           
endmodule            