��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G0��@h ���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����T�l䮱2�W�K��N<��;���Z��4d��{�
��|��Ȋ)zo1���á�x:��*���#�� P���ı���$����1�c/~.)��3\�R�F*}�c}��uOA�ٗ��J��~v��QU���T���딣0&_���X0���2|	p��rw@	@us�犱t��M,�ii^sZ��yq�`݊�|���"rG�
���}�\�.�DV	��dU�;�\�]���џ�_�v%�]��4�:j�l�,9��I{��8�H��s8[Z��pM�i?��n;�|-���g]���͸`q��9`�h[�c�3�n!?0{l�E>�ڹ��o�/*0�(b�شW4;�&�'����d�	�M]�Sw�C/��!��}9���S岦�%I^��������裐d5���Xf/vA�VG��ΊՉ���9?�\�N�{}�=�v��}�����Fz�!�`�(i3!�`�(i3���D��ܒ���-=*�ўo7 ��r曍����&�E����F\F�e���n:�Feb�:8��( O¡0-x����vH<:�wx0�<��W�)��!�`�(i3!�`�(i3�^uf8���m��k��,Ks�k��'?"ӌR�*Zc���6Y��7��8�zv���
����!�`�(i3!�`�(i3�K�Ǔ�\G+���폂P$��j����D��ܒ�cω���s��� ���G����w���*bSl_Ǒ��\�w\_�Z_!1�y~�-�D����K�BB$�W%oY���1:O	��Ѣ�ׇӭ��!�`�(i3!�`�(i3�R�~WI5�z:�ե�F8���m��_g��$o�{V�{��7����6�oр�|D!�`�(i3!�`�(i3�f��mt�5Ә�(�N����4�U]��#��F���j�3����t`�;�rׇӭ��!�`�(i3!�`�(i3����n,��>]��e�?�o�d�I,�D�y:#9�]�B���YH�<,r��,�4�������:�Z����&s�8�e�V�{�������e^KW����Q���D��ܒch?�bnx�˞)��^!�`�(i3!�`�(i3I������e��*�P} ˃$����ܜ?n昼�2#:�ֵ*&E�^8	������hÝ�M���AF�����c��(r6ˈ�z{FQ���'������Fz�!�`�(i3!�`�(i3R�.���2"�k:�Kaw����⤚�[?A�%�Rs{:��r5DE��7a����ZV�o�sȸ�"rR!�`�(i3Ѵ �nӼQ�c�6�fSTK�m�S`j�C��įA��Vq�|`kK��I�t����ۀf|���׎��ax�.Ô�9���v�f]�_�����`���PY�ׯ
`�!�`�(i3!�`�(i3��}2M�; �x����VY7�7Tt��<��d����J�c��ړ!O|V"�����Fz�!�`�(i3!�`�(i3mI��t�����¶o'MrAw&�9˝Sz��E�4.@�����G�������/*0�(b��g��k���M���ʜ�7�]X]���H�B�ׇӭ��!�`�(i3!�`�(i3��_�����v�����������U��5�D�v�l�Ū�TD���	�����v��~��dme����	2�R��y�,��/�􅺊i<�� 7�4�菚![J�i c�i#&\` 1�c�7R/����Fz�!�`�(i3!�`�(i3���KN[tM��.���e�_Mn��"�=��L߇=��ڨ �ߣ�������Fz�!�`�(i3!�`�(i3�(��@'�1����
_cW��jGpș�=���g�H�����tfD?ړ���!�`�(i3!�`�(i3?�k�V�?�����@���#t�Op�ʂ҅��gdjY��<%+�z��4�4���UZ��n9�W�H{�!�`�(i3!�`�(i3��������E����AM��ج��θv���#�%?1���4��%�p�0ΑY3*��K�y؄@�!�`�(i3!�`�(i3�u'JT5��qy�:�ԭsƁ�@����<.���+��T���jB�Fg�Y씤`��px��.��r�M$�*cW)�w�%H�!���Ȗ��h�}�_0+��Zk ��U{����q_H�Э�LP�/�H
M��ވ�c�F�=o����"���	x]̍��;����k�7ꦍzlQXL����g&���ϙc�IK#���{��O��qC*�A�=#+����D�`5�vA�VG��M,������~�*g������_et�rZ�?ђ��P^(����gi���$R���b�>�oa.4��ۙ��x?�s�2zs���T�j�ߣR��zF�Y ��C���!�`�(i3=]A��O�T�`�[�����p:}�L���)	�8V�2�ԧ�fQX��G-�3��rD���Rb��Y�W�7��A�. �*rcxm�N�ɴ��~襊s�� �����p��� [�E� '���I����=��A]�;�J]�r4EG��L����~T�]/L!e*���e��)j��ӌ@�۰V��L { �6��}��%%��c�'GcoTAk�?������F`πѾ��/@��0e��H촼"g&�w)���Hѐ��tAa�/g�P�,-e�]Q��s,�~TM�e�w�G3�E��])v;P���i)���zռ��+��~��'���m�!=�y����h�}
�ԟ�dIQ�0^��-�:L�����Sd,�ϱ���	���Ģ/*0�(bq�� &@RfB�y�I[���b�/'��n9� �1�@tb��?�~���?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�@���rQik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW?���ʢG�M._�I�`D�V�U�'f�ٵ��xMB�9}��DG> �f�������7�����H�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR@�/-��E]o��in�m��+�<4��ˌ�ň��h������R��L�Y�͋�<����d���q����c��� �7ht��}j!�`�(i3���D	��U}c\(�T]�~���nfx�P �ѥ��/�MK�h� )������&!�`�(i3±�sR�{F��JG���%>%��K�h� )g���DD60)���yW�7�ܥ��2�NTګ'6�"dR��|]�������e^KW����Q�E����FQL&�v��H�	A��񊽫wH�HͶ���ܜ?n昼�2#:� ���3�ҺMC�^�.�]`�U+�PA?���\z-��EM���
+����rx�]�V��\#O���o��(�I(�?���\z-ܘ�u}����!�`�(i3x�]�V��\#O���oY{Y����H��c%�ݿ�	�Y��{?a� ~>>ը܅%Gb=]A��O�T�`�[����ЉyE�gr����9�zI�	u)3�!�`�(i3±�sR�{F��JG���%>%��V����D�GX%���d��$���!�±�sR�{F��JG���%>%��������!��B��ҏ�<
DN��b9���A����
��&��3J��\G�Y#�u�'�'�7��r�=�o��C!T*�q���U�ЂDa��(����AA,<��z��}�\w��0]0��l!���?�{�T�	yhPGl݀K�6[��u�(��6���ҋX����>��l%i�-X�Ѕn��ͧ���)�b��|2��w�>8k�(�y��]�!����M[��Ǣ�r����O¶��r�`'���Xw�R� v+0x􈸓��-���{l�f|�ό���.ӽ����
3�i�ҋX����>��l%i�-���E?���Aȧ��b��x����C�*�%.��}���^��W�/��W���5u���贕ƫ�ܶ	´@x�p�M@�� *����{l�f|��rs�i�/ �m^'����ܜ?n昼�2#:�G�&�;?�Q^�MY:+:  E��a(􆿳�ؖ��d�I�� �:&�����ˉ�1�:�Ω�s8�R�	�}����T�l䮱2�W�K����Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�$:v��`E�EYZ/�h�@�o��I�?g�f���\X�<����8��U�[��Egܹ���fq�Sy�������Q����H	+��j��B�v�(Ȣ4 u�>�QB�{\��Q�U�;� *ӄhE`Ԏ��%�R�C�'f�R6�1����י�L����-�8�X���開#c���܎��/!Di�����+�� �q7�F ��W�A#Yl6���@��+Te�vWi���������5	��)��8'V����(��1੡�3����Β �GG�7�)��5����`K_T���0��x�]�V�����ɢݣ2l|�*"k���(ӈ��Q'�y>�1!������d`O��� ��b�FP&(����/�7�d�٣��c�A�L'�}g6��g���cH����\�悽I��y��,H/�� ��b�FP&�%5:�����d�٣��c�A�L'�}g6��g�Njn����yO�E���%�;���EWr��U�L��Z��cfo�w��.�`��+x�r���?���������OZ鎬�������(�����K�J��8&���I���8|�W��{q3�e�[=F���-/a8[��p#ِ.�����	����@|����r�����\}{���b�/�J�mx޴,��$e�z8_��ݚ�Н�����$K7͍��B0�����V�;b�-�2�'{w#/ B�@�І�y��ˇ�h�����?S�� #�K�DQ�����M��%�p@<�6�Q=��� ��RiS@���;b�-�2��;�P�t�5�W�fD��0��ϼ%�bu7���Q�s�rs�i�Zy�ҠE�W5_�D8��SENan&��u�Y�KG���;���o*A&-�Ri�5����f���s,�f��b~�]S�8=��䅿��nz[�چ�v�9��8�w��U�%D�)&���ݚ�Н�(*�O�qܴr���[}�N�`2���K����b+}y[!�`�(i3��!�����&~e�e��E{��hC>���d���|e"ʁ���MյxZ�6��	Ղ�I8�y\��S��z��Q���!�`�(i3U /숇�v-�^�L�-�;S5b	��T�.����j��6����&kQ�fY�U젩`#FW8�	��PGc��WI��}Dq�f�G�&ց�*�ny/f!�in���}���S.�3����7�!C�!�`�(i3pı��0����{%F�Z��3��w��\�Wݺ���� f�ݓ�W���,�GV��4�0 L?ஹ�%��\,!` 5(��ݚ�Н�(*�O�q�b:�<�ۯ�[}�N�`2���K��h��'���!�`�(i3Gٙ�;y��&~e�e��E{��h�Oz5@p~���|e"ʁ���MյJ�h$"h>�	Ղ�I8�y\��S��z��s���
��!�`�(i3U /숇̷�%�:�-�;S5b	��T�.ęj�+�BU��6��c]Ip���U젩`#FW8�	��uq�B�%���}Dq�f�G�&ց�*�0{�,A~n���}���S.�3���+o��vHm!�`�(i3pı��0���nK�3Z��Z��3��w��\�W�1h��d0y�ݓ�W���U�2<4�0 L?ஹ�%��KvfЗ��ݚ�Н�(*�O�q1��h��ˀ[}�N�`2���K��g�6~x��!�`�(i3� ��F�fM&2A;~N�E{��h1�����
���|e"����1��eǡ��=ֺ��W0�]��x@���37y����m�/
?�E�i�m}6O�D mWNTT7���1�a�;q(�I8�G-��)IMdK�Ch���UJZW��sT��E����F�t�t>
x�Pumi��|���jL#{��X:g��}�
�?���l�(�2#��4r<{������3ό���.���g�,P�nw�����A�?���0yV�6IWJE�!r}<ﷹ�t�Z�f����@1��?�T�\ �ͻIb����rs�i�/ �m^'��D24N<I8����\.W^�V]��}R�wX��}�
�?�套�qD0���HՕ�O�M:R	�'����Ԝ��I���X������@�&_E�EYZ/���V�	�Ncny��&�;a"��0�혅vº��żפ	�?9Pjp��17e��:r����ZqJ?�d���&��ꢤ�Og1����?���zf�l�=_�#<����k�5,���������9b�S� 7�v�ԯȥ�����S�7>�����ǚr��yݒ'��Ң>AV��	��y ��f"�:�HCaIMlP.s~#hdbO¯Fs̃\��W����2D)ĞSy7[��7%^�,ף썚vյ[+8�G*8� �k����#M/�����.�̓l*>+6�����C#/<���qk˹@��]&�2�Ɏj���|��p?�yG�<Y���m�F��?3�t6��y�~?�2vŀ�#����zl��U�2X���#H�S��mr>���*��~E�_�#<���ӟ@^9�C�Q��JsyLJ��=?*럐D�f�.��^j��R��(%�2Y4M��U��)���Y;e�iK-pm!9�>��`UNP��q��É~�nJb�G �!�`�(i3$�xKw�6��/B����~?H�?�����3@�4��r:O��%(���1�'�p[�8���&��~�26��\2|Oo�{b�!�`�(i3��os�z���}Dq�f� ��b�FP&t�G���f70����a�\����N'�D��غ���"��~�26��\\��;/���*e>�{,ԯ���gnņ��#�b���$�Qu�R�47��vL n9-�Nû9Z!�7U��sB��򨂓�m@Ǒ�5�o��7��E����F����o<rS�b�8Z���oگ��r���%��Q^�MY:��H<㕕ѿK��#�$����v�B���(�_���ߦ�D��.�E����F[s�9�-n���~�2�?�B�����lC��U�T�\ ���:5A��p�~�26��\����g"m�	ǰ�O�l�7#.�KUfc�^�X�{��=��$�Qu�(N��LI��$"�(z�J��Ҕ��i�ϕ�"��,۽��������y�(����<m�df�L�_dj�Ï��	�l�lM�3 H�RtV�^v�t�J��0s�J(|&�@Sހ#��_H�RtV�^a3@��[/�L��O��p�`��q�':E��nd_�oD�a���裣2�`r-��&�X�P�|��]6���k�T�A�}f�֠�e�ޔ*����!F�G�`���S����\e&���m�?�϶q�U��!�`�(i3�i7N�_�wDo�h�'�t�Z�f�t���p,�7�g��U-�egt�n���!�`�(i3���F1������$����iVMՈA��'''���:�JK�K�r��Lm�:�w��Ip�
�:qEpCt�w#��@�ݚ�Н����F1��kټ�b�	�RCJ�����@�ĵm�ݚ�Н����F1���Q����>��&#��B�[�g�DPp�HN��R��bP�63Z�tp�8��7���@�e
@t�G�����,1�!�`�(i3U�	Y���a3@��[/�L��O��p|���_��}["��4��:��Kd�CN�zB����Ȋ�?ӳ4�;Ⓠޕ;j�j�������"�
�T�r�5��� л���}��!�`�(i3�JO�'��+��K�L�Ik�GIJ�,��=��i!�`�(i3�JO�'��`gw�T�с֜>�E�2w�f�%!�`�(i3<p,�mY!q�`�	6�����Ȋ�?ӳ4�;Ⓠ�X/�7�D(hþ�f�<z����Uv~��6������S>�y�-�RJ5Y�bv�N�ԑP�מ�����y��lD�f=R����X������%A,�ι�S�t)��:5A��p�Y(��<��4�;Ⓠޕ;j�j�������"�
�T�r�5��� л��r����0�	�:]I1}�ั):9��tf��!���i��L��?����9��v�9��a3@��[/�L��O��p��?z��t�g"m�	�uE9�+�廻��j����Z�!���6������S>�;�u��tF�{F#��~�>�R�����6������S>�y�-�RJ5Y�bv�N�ԑP�מ�����y��lD�NA�1;S����Yk��1}�ั):9��tf��!���i��L���2���l���}Dq�f�1}�ั):9��tf��!��Ϗ�2�ed4���Ȝ�}Dq�f����E?��1�a�J������;c�~��=�g�żפ	�?9Pjp������PN��7�v�ԯA��bu�x��ݚ�Н�S/���]˝Sz��E�4.@��:u]R��GX�Z�X�W�NY���eb��D@f򨞊i���)=�,J�� ��C���򨞊i�����-����!�`�(i3ˣa7κ=�c�W���c�/_����^�'�)�Բc1����?��S(�`�ՙ!�`�(i3���F1������$��\R�j°��ݚ�Н��̢k���!r}<ﷹ�Q^�MY:T1�Ɓj9��jg����ΒՎ h.\���Z�
,�/>��a���9w��d���[�,�/>��a�r���m�5��ݚ�Н� As�Uq	�*��D�x�Ěο��h�SJr~�PQ%cp��g��v�9��!�`�(i3�JO�'��qc�Vۍ�پ�[�_��!�`�(i3����١�$�ݛ5�CNi~�N,7tL���4X%��C_=A�H�RtV�^����&��vL n9-�N*��D�x���Q���kO��u�:�HCaIMl�i;��B��}Dq�f�`
 ֢��؜J��v,ŋ�����)�W�=�k��:5A��p�Ra])n#����m?�V?��?s��Ԏ����:v~E�)d,%B�����ݚ�Н�h큈���g�W����w:�눔�C.�u�X��I�ՠ��t����>PQ%cp��g�H���~��!�`�(i3E��\�����7}#�ouߗN���g�3$�J�5'!�`�(i3��Ě�����}Dq�f�a3@��[/�L��O��p��?z��t�g"m�	�uE9�+��HN��R��Gu�"�0�`
 ֢��)�at��*��;@�1��/}�׏)#uE9�+����Ě����E�i�m}6߸��S�Ȍi��(.�j2����j�F8aT��3G?�d���&�bO¯Fs̼�v��z�=�v�U�φ��<�6�$>ʹ�*�Ĺk\������`�5Ԍ������E����Fxy0�u��¤M�[�g��DW��ԅ1Qr��[��l_ ��b�FP&p�]f�"v!�`�(i3���7���~ֱ�q�����2�w�] O�m�;�ٜ��׽X���K�J���N}�m��{W`�v�L���f70���i3<�f�D.`�Z���N}�m��{sy�,"��f70���i3<�f�D.`�Z���N}�m��{ڃj��-��\����i3<�f�D.`�Z���N}�m��{��{&<c�yQ���4�l��qBVF��`���oN}�m��{zh��ʊw!�`�(i3=]A��O�T8�G��oBߓ��A}:h:
���9
!�˝Sz��E�4.@�o-�!���H�g��U-�e��,H/�� ��b�FP&]���6d�!�`�(i3�I��?��\/ �m^'��D24N<I8����\.W��"X��[��Q[R�7N}�m��{n&��Y����o�x���i3<�f�D5��E	c�H�\��;�,�~�26��\��r����g"m�	ǰ�O�l�7#.�KUfc�^�cQ�0.��èVe�;ed ̅��Ȝx�5W ��̫(� h�ҩ�|��^���#hM�\���|��^���#�� MQ�S>������:
��x�{�\��N�Ś�-����;�jmT�#3M)Q;�.��1�{��(���XW�G�<I/��\]� h�ҩεSENan&���ߊ�ֲ���ܜ?n昼�2#:�^�V]��}>�C�;�����:=����l��+� �z����	2�R�(�p���&l�b�u�!�`�(i3�������l�����)l��4���O�>�k}�r��N����󑩄�n,��>]��eW���ђ״�~�YI�!�`�(i3�m����9N���{��c����'�u�
rx�pj�d!�`�(i3���Ȋ�?ӳ4�;Ⓠ�:�7jZ[r�.-�gg$Zzr�!Xk(��A,Q�mr�ݚ�Н���6������S>���S��a�bv�N�ԑP�מ��!�`�(i3$f��_Ub�F�S�1 �����l������6z:�B����]��V����l���.�et�rZ�?ђ��P^(�՘�}���������J�\���=��}���)��U�UH�RtV�^!�`�(i3z���r#� ?����6	�T��u~��t����>PQ%cp��g�H���~��!�`�(i3���F1������$��\R�j°��ݚ�Н��Ra])n#����0�������ߺ��8�ۦ�P�X��P�������pC-��h�>
A��%���'��eEqWU���>
A��%��WG���;� h�ҩ�!�`�(i3k�s�X�C�GM��4�ūd���8tO�M:R	�@tqx���!�`�(i3`
 ֢��؜J��v�S1��6�uE9�+��!�`�(i3����١�$�ݛ5�CNi~�N,7tL���4X%��C_=A�H�RtV�^!�`�(i3
Cj�R[z�(�� '�i�*ڃ݂S�����3�t�.K��ߎ�x��y��v�9��!�`�(i31}�ั):9��tf��!
Cj�R[z�!�`_q�!�`�(i3�̢k����J�\���=��}���*rcxm�N�e�{�W!�`�(i3h큈���g�W����w:�눔�C.�u�X��I�ՠ��t����>PQ%cp��g�H���~��!�`�(i3���F1������$��P"G�wk��=MNԅ,+��}Dq�f����%>�rGO�D mWN!�`�(i3��֖+�){?a� ~>>ը܅%GbNÌ�Y,�u��r��!�`�(i31٥xu5=�Р��U�1Q�\��^����!�`�(i3�	��x��ݚ�Н�����l�鉌(*$ΐI�q����!�`�(i3c���P�vћv\���7��{����S����9�@��!�`�(i3`
 ֢��؜J��vv��v�K���x����VY�l��NI��ݚ�Н�
�:qEp�;�P�t�5!�`�(i3$f��_Ub�F�S�1 �fĉ>99��R�Q���~��p�������l���7�����Vq�|`kK��I� zSd��;��-����!�`�(i31٥xu5=�Р��U�1Q�\��^����!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ6�v�Lv v|��V��*�R�~WI5�T�ϓ9��IX0F�MV�ҁGG�K�BN
\��=2�L-�f���f\�i��W�x]��0�N}�m��{W`�v�L���	�zQ�$Y	�I]����2N��n�ܖ �&���J�p��2,��T���$�Qu�Y��m���Y�B�N�����wRy�����q8n(�E�K�.�O��_�8&���I��S�J\7�_�Ƭ7~��J��V�ShT������qD��=a�^7�1tSjv�N������{��7�f�8
��u��r���n��Nh�^"�Y�.����n�f���fv�$� ��n=n�k-�;��H`��!�οn>a3�qj&�G�;�jmT�#�&5�/h/�[�a��O��_��-����!�`�(i3f퀔����W����Qy +߂X}����eՍ�s�)\��w���f\P�.��$�'�ͬ���~,�H�͛����%>�rGO�D mWNHN��R��bP�63Z�t����g�Z��3��a���!@�f")u��r���9�Uv~'қ�-��F4��5�\"^�� h�ҩζ
�t��T&��ۥ`�M?��y�!�`�(i3�U�{��YD�íN=]b~*��s���?����2vr5�Dѯ��B� �b��!�`�(i3<���K<�Vq�|`kK��I����<����1tSjv�!�`�(i3� ͷ�	�������e�؟�r���������+ot����m�����r����!�`�(i3�R'cf��i�X!�!D��(J�f�x��2�+�T�\ ��[��(��!�`�(i3�y��j��k�=��7���P%�H��Jq��BѲ�+���L>!�`�(i3��6��w=\��*ȜD���|�]�)�Z����J�]�]K����J��!�`�(i3!�`�(i33���Z��$����꨽X�4�M���)/��:5A��p!�`�(i3���W0�]��x@��!�`�(i3.��J�޺��:p~	E�<l��uE9�+��!�`�(i3�d��R�;Fc/�p@�dB<4RW��rS�b�8Z��W�6?��O�M:R	���;Opr!�`�(i3!�`�(i3M���CO|e��߬/�~8���|A�W'
SxtC��)� I��r��P��ap�7?�A���.��r�ݳ�sO�~�fBǂ<�'�/��YF�"�߼����(�%���]v1�_ُE2�DZ��DO��"hń��0͕s�i��\����4q�.-�gg$e���K��!LtD9$Ο�
��[H~����}Dq�f�!�`�(i3fF�5.]����C�i��^!�`�(i3�	��x��ݚ�Н����y��lDlڍ��p�|92w$�P3z}�&�!�`�(i33���Z��$����꨽X�4�M���)/��:5A��p!�`�(i35���eH��_
�5Y9^��
Li�#fC�V��a;����Yk��!�`�(i33���Z��$����꨽X�4�M���)/��:5A��p!�`�(i3�?�JY�)�q��ڍ!�`�(i3�i7N�_�wDo�h�'�t�Z�f�t���p,�7�g��U-�egt�n���!�`�(i3�/��@����*��Sx֐�M�4m��?�N����!�`�(i3�'ѧۂ��#����E������C.�uE���h�/	��26h�W�5��|�F��|�'�&|e��߬/�~8���|A�W'
SxtC��)� I��r��P��ap�7?�A���.��r�ݳ�sO�~�fBǂ<�'�/��YF�"�߼����(�%���]v1�_ُE2�DZ��DO��"hń��0͕s�i��\����4q�.-�gg$e���K��!LtD9$Ο�
��[H~����}Dq�f�!�`�(i3fF�5.]����C�i��^!�`�(i3HN��R��bP�63Z�t���%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��j�_�Ƭ7~��J��V��L֞S���`����ǆ| c�]hgi�K�%@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���j
�D