��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G0��@h ���iQ�����-v�ZN��p]e�km?Ix�J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lV�t�[;�Z��4d���Ġ���딣0&_���X0���2|	p��rw@	@us�犱t��M,�ii^sZ��yq�`݊�|���"rG�
���}�\�.�DV	��dU�;�\��I��Sf	��,h;2���۟�
$�e
�9��Ax!P����9SA���S�BgV�0�ם�kk���6 xI+r�� 0�D�A�f�mX��)D�b@���R��c��@0����{K��"\��7B ��IB~���P���	Oe�P(�[/ C]$�%{��N3y��	8��i�xx�j�GEc�0��˩���.|�-J(��6�&�]���@�3�gĸ����P=�%u�:��\[�K����T�F�8t$/�:M7bR�&	��/v��~38C�	��x<�Ⱖ�(��.2�@���'�.���1Ԕy\ �პ��K��Q�Y�:��.�>r7��oݮC^eG=C�T��4�����uS�+].�/��	c��Y�sVh�a�ei�P�?�_��,���4�8t��^�?!�ܵ�c8)9��?{�5�V���W���/����Ӊ>H0�^Лq>�H6�կ��xju�^u�b�`$�Ƣ�/��_a;�+kB�����H&���@�>� ��o����;%�1��wd7>Q�U��y�@{���g��Q0�@���rah�oY���3��DX�\7Q��^�Kp�?����&ʇ�k2(
����R�g#��������UE�R�D[�?�٥�ٽ�@�������ꏶ�=��g���g����+ ���r� �'�f�!�@ٰ�Ř�h^����y�	W�%N�=�Db妘jC�
����١�=FRѼ���8Cv�c
�������K��S�����a�7�I�E�-�iׂ�r}�̤뢲�
�A��߱��Wf'�j�"�r�47�p��M�VB�p���[�1T{pў�%63T�N�+[�����,[$~������ �Nb)�w�od[?�j���+�x�K�#��m����7ɥ�׋�ޒ}12�}��ɣn�Tn���i�i՞Q�o�~����p��_Q�!�o_�SW<*
0���ۭ�
ۂ>F�%}/h-��]m���/�9ӯ�1�(1�Y�9J��Iǋ�Oi-*���i <��Mr�J�M�D�9Tp��C��u�9"5�$9XK��w�\�\��M�������m�����,o
���開xm��D�褐�2��ql5���erK�^��l�[//Vq�|���۶+M��Gq*�r�c�y���X׼p�Nģ�Z�8��D���pߣ��G���a����	�y{y�Zw�E�!��,h;��}	�l*Y���KS�p\�5K���6�� "Z����.���\��Wg֘m��R�G�)q@�Wԏ�6{5-Q��]����>�LT<��k2(
��yTœ�(]��,sȸ�"rRZ���@��E� �/�z�
>�"S@�"� �K� w�;�d���N�tכ݁=9�|Z���ߐ'�[�Z���1VU���+L��h��X�vB#|y{����P7�.yt�gU*Z9B[�^������+�ͫUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�#CC1X�G�ۄ��O���azhݪm����Y�{'%s#K�v]|nf<�,=K�F��N��j��D���s���ئS��.V&��B֥�(����5��M�=��S�=hd��1}Kط��4q������Tkd�_���n���	h��IB��XP���<����k�|�c8?-+eN7��c��;��\�vŮ�@W��C#/<���q�V�&��'�E����#3Y��P4p�ji�ШFs��X�vHޓh`����W�3�~�B�6��J���Z/���V�/��M?� g0/p�i�F�s�3�̞~%������a[�x�۶�kvɎ����9-�8���� �@��&}"	�c�o|e.��xu	���S8�
T�F�����lC��U�T�\ ���A����l��4:�CTv�ј�"��Z鎬�������(���/p���x�CyW�f�tR�wX��DsQ�V�r[1B�VtE�<��z��}�\w��0]Y��
�iC�E����F��j��\w��0]%��C���+�
�c�~��j��\w��0]��0�&�ͭ�E����F��j��\w��0]{k�h�+m��q'��7G#+�Ǘ0z�cUL
 '&1���D���J��8���/��-�
�]o��in�m��+�ވΦ�籢ֺ�9H��/ Oag���:tӫ�C+��T���.��Б����K��!Z�NCIw4�dט�w���۴��pD��/��+JHn��z�'8^�#ٸ�U��֜��3��pKU��G��{Ǧ%W& s���r7�����^���I�� ��˽��r��B������8X�ŵ���XP���rS�b�8Z���'�e�����"�?;(��j67� ��˽��r��B�����)c��jCIÙ=�H60���	��p�(�oE��(��f��Q�m��'A>\^M�Ɣ�5����`K�������$��\�v�n��j�S��(��ir������y�$�g?_��<'P��!jcCA�T�g�v�'s��k� r7�r��#[^]�Z����Pcsù�Ln��S�WHWG��i�IW& s���J>:F5q�E�_s��G�b!��u�!-B=�6f5בvk!7s�9���o��S8�9���SN��'6���;8=�g��U-�e,%�0g���[�=�5x���?!6)X��-�>�Z鎬�������(������oD��;mQ��8���/����,DpR���ע�!OF����+�J��Y�{'%s�rOw���é#7ۏs|�L;Л��|#9���b!��u፬!#��Rh�\�٬y�7s�9���o��S8�.�9�T�����k��$a(􆿳���2����..W���ۗACd�\��"�,�>E���]�!��	Ǹ�y85�2�N�Wb�2��Я�R�wX��}�
�?�<��0n|�!h�b���t��!�=6s{�0z�cULn�4Z_U���l����g��U-�e,%�0g���l������*b��93�|q��-��Z鎬�������(������oD2��Я�R�wX�չo��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�_-�B'�b�@�|�S��*��B?���4U1������E1�y�WQ��KF9q��>j��(���ll�!(�ʕEr5��Kr���N����+Ed�J�5����d�φ_i�����؈J_�P��ዧ3��^�y�b�5�!�� %	���{ s�3*(�{�DPx�V���R��)�ޔ@��|��:`2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���X`
�t%>^�ߒ.�qO���WS���
���A����|�������-�YM*b��93��bj����kѶ���� >�������.�Ӂv��9Kd��"�����ڗ�\���V2���<�؊�"�Dz�Q��y{y����x��F�U| c�]h�G2[�4��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��.2�@��Me�A��.X���Y �?���M��,:�-���F����D���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�0�"�!S�ff�݃v{��lw	V��aD"�'6���;8=�g��U-�eӢl*H0*�T�'Y�����ⓚ��ToME1�Pcsù�NdE��Q���;mQ��b�c��=9�ߨ�,R�e>۵��>�}�r�KņMC@����^�	I�����k��$a(􆿳�eJ�Í6�U�N��S�Ԍ��e�[�0v��t���1�����ׂ�⾉�ƃ
ᾆ�x�S�v�b�k�#7ۏs|�:�9,�52�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ���q)2���8
[#oAp)U��zN���]$�%{[�a�(�����9��J�Iܤ�����o�5�;2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�^�wo���Z��	�`DÜk�K��h̷_��yC��S8�\�w�4�*)�2�"ղ]�6��2�~�P��qa���=7�;-�]����2jɸ�2�V��ᄲ-��B?-XK���jVѭ@!�`�(i3!�`�(i3�ui|Ɏ;�0z�cUL��ddՅ<Ta��;���=�[%�('T����7 �>N��bz�9ڈ�KK?B�5 �8��B��j	WJ�u���������-��d�H�����'���Xw�j�7��AԢ�a\�#P��W��������|Pcsù�u�ȭ�>�W��7(�bOh[X܉]�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�a�}�$��W�6?���N��S��pP�Fc�����k��$�����k�A#�G=�]Y�����Y&X?r>幛o1����k$ !�`�(i3!�`�(i3�]�!��	Ǹ�y85��X��I�ՠ���aٔ^?��[+��.Ȉ�;1�˚�!��JlR�`<Y��sp@�9�m{�L�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3AԢ�a\����R�?�������|Pcsù�u�ȭ�>ѯN��S����%����<��0n|�!h�b���t�j��s/�rs�i� S�xSVe�W�6?��W��7(�bOpP�Fc�����k��$����导�?!6)X�Yկ����!�`�(i3!�`�(i3!�`�(i3!�`�(i36�&��=�'�)�Բck�A#�G=���%A������D�ϲ]�6��2g�1�9�UkQ���7�!�`�(i3!�`�(i3!�`�(i3!�`�(i3k,q�*��	���3\�a%,ʋ�j���jVѭ@!�`�(i3!�`�(i3�ui|Ɏ;�0z�cUL��ddՅ<T]v1�_ُ�T�'Y��Y��{&���'6���;8=� ��g�SEս�9�j�x*�����!�`�(i3!�`�(i3!�`�(i3!�`�(i3�uz�#-]iL�1p/-�����̵?o����oD�d5z�R��5 �8��B��B�n��َm(5!�`�(i3!�`�(i3!�`�(i3!�`�(i3́1)�V9�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �����:8E��)$F"�h\A�/�*����7/���mX�T�h��ϾL8��}��ɣ����0��B��!1n�r�9e���ƽ>j�(d:Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�#~.��,�IX0F�M�U��)���Y;e�iKI/B޾Pb�i0[���S�J\7&���"�g7w?��|����gmJ/���'ž1�|�'����z.��W��!�`�(i3����j��3���B[=����e���A��s�R�b>3��g�2��}��D�o�&x����E2b�z'hۉ)��d�7�q��k��^�1��dc�@c�����h�'�ɳ��<�6�Q=��ž�Ć�T���7X���c�}�:
��x�{�\��N�Ś�-����;�jmT�#<��0n|�!y6]�o���s L�Zl�WG��Hb� h�ҩ�?V��j�c]���I���������h)C!nk��q-K���չ�>ʰ��ߨ�,R���"X��[��Q[R�7՝� s�#���k$ ?V��j�c]���I���������h)R�Rl��K���չ�>ʰ��ߨ�,R���"X��[��Q[R�7���%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��j&���"�g7w?��|���.߅�[j'�_2��VU(��z�j�6f�L��.